Current Comparator Simulation
* this file edited to remove everything not in tt lib
* .lib "./sky130_fd_pr/models/sky130.lib.spice" tt
.lib "/Users/rej/.volare/sky130A/libs.tech/ngspice/sky130.lib.spice" tt

* instantiate the Current Comparator
Xcmp Out X0 X1 X2 X3 X4 X5 X6 X7 Y0 Y1 Y2 Y3 Y4 Y5 Y6 Y7 OutCmp InCmp VGND VPWR tt_um_rejunity_current_cmp

.subckt tt_um_rejunity_current_cmp ua[0] uio_in[7] uio_in[6] uio_in[5] uio_in[4] uio_in[3] uio_in[2] uio_in[1] uio_in[0] ui_in[7] ui_in[6] ui_in[5] ui_in[4] ui_in[3] ui_in[2] ui_in[1] ui_in[0] ua[2] ua[3] VGND VPWR

* NGSPICE file created from tt_um_rejunity_current_cmp.ext - technology: sky130A

X0 a_21880_41750# a_21880_41750# VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.35 pd=2.7 as=0.4 ps=2.8 w=1 l=0.15
X1 a_21880_41750# a_22050_39050# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.54 as=0.168 ps=1.64 w=0.42 l=0.15
R0 uio_in[0] a_23490_39050# sky130_fd_pr__res_generic_m2 w=0.45 l=0.05
X2 a_21880_41750# a_22530_39050# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.54 as=0.168 ps=1.64 w=0.42 l=0.15
X3 a_24200_41490# a_24200_41490# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.54 as=0.168 ps=1.64 w=0.42 l=0.15
X4 a_21880_39160# a_21880_39160# VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.35 pd=2.7 as=0.4 ps=2.8 w=1 l=0.15
X5 a_21880_39160# a_22050_39050# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.54 as=0.168 ps=1.64 w=0.42 l=0.15
X6 a_21880_39160# a_21880_39160# VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.35 pd=2.7 as=0.4 ps=2.8 w=1 l=0.15
X7 a_24200_38900# a_25610_39160# VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.35 pd=2.7 as=0.4 ps=2.8 w=1 l=0.15
X8 a_21880_39160# a_22530_39050# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.54 as=0.168 ps=1.64 w=0.42 l=0.15
X9 a_24200_38900# a_24200_38900# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.54 as=0.168 ps=1.64 w=0.42 l=0.15
X10 a_24200_41490# a_25370_39160# VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.35 pd=2.7 as=0.4 ps=2.8 w=1 l=0.15
X11 a_23810_40680# ua[1] VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.45 pd=2.9 as=0.4 ps=2.8 w=1 l=0.15
X12 ua[3] a_21570_2680# VGND VPWR sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.8 ps=3.6 w=1 l=0.15
X13 a_24200_41490# a_25850_39160# VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.35 pd=2.7 as=0.4 ps=2.8 w=1 l=0.15
X14 a_24200_41490# a_24410_39160# VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.35 pd=2.7 as=0.4 ps=2.8 w=1 l=0.15
X15 a_24200_41490# a_24200_41490# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.54 as=0.168 ps=1.64 w=0.42 l=0.15
X16 a_23810_40680# ua[1] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.189 pd=1.74 as=0.168 ps=1.64 w=0.42 l=0.15
X17 a_24200_41490# a_24890_39160# VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.35 pd=2.7 as=0.4 ps=2.8 w=1 l=0.15
X18 a_24200_41490# a_24200_41490# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.54 as=0.168 ps=1.64 w=0.42 l=0.15
X19 a_24200_41490# a_24200_41490# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.54 as=0.168 ps=1.64 w=0.42 l=0.15
X20 a_24200_38900# a_25370_39160# VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.35 pd=2.7 as=0.4 ps=2.8 w=1 l=0.15
X21 a_24200_38900# a_24200_38900# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.54 as=0.168 ps=1.64 w=0.42 l=0.15
X22 ua[3] a_21570_2680# VPWR VGND sky130_fd_pr__nfet_01v8 ad=0.168 pd=1.64 as=0.189 ps=1.74 w=0.42 l=0.15
R1 uio_in[5] a_22290_39050# sky130_fd_pr__res_generic_m2 w=0.45 l=0.05
X23 a_24200_41490# a_24200_41490# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.54 as=0.168 ps=1.64 w=0.42 l=0.15
X24 ua[1] a_23810_40680# VGND VPWR sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.8 ps=3.6 w=1 l=0.15
X25 a_24200_38900# a_25850_39160# VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.35 pd=2.7 as=0.4 ps=2.8 w=1 l=0.15
X26 a_24200_38900# a_24200_38900# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.54 as=0.168 ps=1.64 w=0.42 l=0.15
X27 a_24200_38900# a_24200_38900# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.54 as=0.168 ps=1.64 w=0.42 l=0.15
X28 a_21570_2680# ua[3] VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.45 pd=2.9 as=0.4 ps=2.8 w=1 l=0.15
X29 a_24200_41490# a_25130_39160# VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.35 pd=2.7 as=0.4 ps=2.8 w=1 l=0.15
X30 a_24200_38900# a_24410_39160# VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.35 pd=2.7 as=0.4 ps=2.8 w=1 l=0.15
X31 a_24200_38900# a_24200_38900# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.54 as=0.168 ps=1.64 w=0.42 l=0.15
X32 ua[1] a_23810_40680# VPWR VGND sky130_fd_pr__nfet_01v8 ad=0.168 pd=1.64 as=0.189 ps=1.74 w=0.42 l=0.15
X33 a_24200_38900# a_24890_39160# VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.35 pd=2.7 as=0.4 ps=2.8 w=1 l=0.15
X34 ua[2] a_21570_2680# VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.45 pd=2.9 as=0.4 ps=2.8 w=1 l=0.15
X35 VGND a_24200_41490# ua[1] VGND sky130_fd_pr__nfet_01v8 ad=0.231 pd=1.94 as=0.231 ps=1.94 w=0.42 l=0.15
X36 a_24200_41490# a_24200_41490# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.54 as=0.168 ps=1.64 w=0.42 l=0.15
X37 a_21570_2680# ua[3] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.189 pd=1.74 as=0.168 ps=1.64 w=0.42 l=0.15
X38 a_24200_41490# a_24650_39160# VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.35 pd=2.7 as=0.4 ps=2.8 w=1 l=0.15
X39 a_24200_38900# a_25130_39160# VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.35 pd=2.7 as=0.4 ps=2.8 w=1 l=0.15
X40 VGND a_24200_38900# ua[1] VGND sky130_fd_pr__nfet_01v8 ad=0.231 pd=1.94 as=0.231 ps=1.94 w=0.42 l=0.15
X41 a_24200_38900# a_24200_38900# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.54 as=0.168 ps=1.64 w=0.42 l=0.15
X42 ua[2] a_21570_2680# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.189 pd=1.74 as=0.168 ps=1.64 w=0.42 l=0.15
X43 a_24200_41490# a_24200_41490# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.54 as=0.168 ps=1.64 w=0.42 l=0.15
X44 a_24200_38900# a_24650_39160# VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.35 pd=2.7 as=0.4 ps=2.8 w=1 l=0.15
X45 a_24200_38900# a_24200_38900# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.54 as=0.168 ps=1.64 w=0.42 l=0.15
R2 uio_in[2] a_23010_39050# sky130_fd_pr__res_generic_m2 w=0.45 l=0.05
R3 ui_in[2] a_25610_39160# sky130_fd_pr__res_generic_m2 w=0.45 l=0.05
R4 ui_in[6] a_24650_39160# sky130_fd_pr__res_generic_m2 w=0.45 l=0.05
X46 a_21880_41750# a_21880_41750# VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.35 pd=2.7 as=0.4 ps=2.8 w=1 l=0.15
X47 a_21880_41750# a_21880_41750# VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.35 pd=2.7 as=0.4 ps=2.8 w=1 l=0.15
R5 ui_in[3] a_25370_39160# sky130_fd_pr__res_generic_m2 w=0.45 l=0.05
X48 a_21880_41750# a_23010_39050# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.54 as=0.168 ps=1.64 w=0.42 l=0.15
R6 ui_in[7] a_24410_39160# sky130_fd_pr__res_generic_m2 w=0.45 l=0.05
X49 a_21880_41750# a_23490_39050# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.54 as=0.168 ps=1.64 w=0.42 l=0.15
X50 a_21880_39160# a_21880_39160# VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.35 pd=2.7 as=0.4 ps=2.8 w=1 l=0.15
X51 a_21880_39160# a_23010_39050# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.54 as=0.168 ps=1.64 w=0.42 l=0.15
R7 uio_in[3] a_22770_39050# sky130_fd_pr__res_generic_m2 w=0.45 l=0.05
X52 a_21880_39160# a_21880_39160# VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.35 pd=2.7 as=0.4 ps=2.8 w=1 l=0.15
X53 a_21880_39160# a_23490_39050# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.54 as=0.168 ps=1.64 w=0.42 l=0.15
R8 uio_in[4] a_22530_39050# sky130_fd_pr__res_generic_m2 w=0.45 l=0.05
X54 a_21880_41750# a_21880_41750# VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.35 pd=2.7 as=0.4 ps=2.8 w=1 l=0.15
X55 a_21880_41750# a_23250_39050# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.54 as=0.168 ps=1.64 w=0.42 l=0.15
R9 ui_in[4] a_25130_39160# sky130_fd_pr__res_generic_m2 w=0.45 l=0.05
R10 ui_in[0] a_26090_39160# sky130_fd_pr__res_generic_m2 w=0.45 l=0.05
X56 a_21880_41750# a_21880_41750# VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.35 pd=2.7 as=0.4 ps=2.8 w=1 l=0.15
X57 ua[0] a_23810_40680# VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.45 pd=2.9 as=0.4 ps=2.8 w=1 l=0.15
X58 a_21880_41750# a_21880_41750# VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.35 pd=2.7 as=0.4 ps=2.8 w=1 l=0.15
X59 ua[1] a_21880_41750# VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.55 pd=3.1 as=0.55 ps=3.1 w=1 l=0.15
X60 a_21880_41750# a_22290_39050# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.54 as=0.168 ps=1.64 w=0.42 l=0.15
X61 a_21880_39160# a_21880_39160# VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.35 pd=2.7 as=0.4 ps=2.8 w=1 l=0.15
X62 a_21880_39160# a_23250_39050# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.54 as=0.168 ps=1.64 w=0.42 l=0.15
X63 a_21880_41750# a_21880_41750# VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.35 pd=2.7 as=0.4 ps=2.8 w=1 l=0.15
X64 a_21880_41750# a_22770_39050# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.54 as=0.168 ps=1.64 w=0.42 l=0.15
X65 a_21880_39160# a_21880_39160# VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.35 pd=2.7 as=0.4 ps=2.8 w=1 l=0.15
X66 a_21880_39160# a_22290_39050# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.54 as=0.168 ps=1.64 w=0.42 l=0.15
R11 uio_in[6] a_22050_39050# sky130_fd_pr__res_generic_m2 w=0.45 l=0.05
R12 ui_in[5] a_24890_39160# sky130_fd_pr__res_generic_m2 w=0.45 l=0.05
X67 a_24200_41490# a_26090_39160# VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.35 pd=2.7 as=0.4 ps=2.8 w=1 l=0.15
X68 ua[0] a_23810_40680# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.189 pd=1.74 as=0.168 ps=1.64 w=0.42 l=0.15
X69 a_21880_39160# a_21880_39160# VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.35 pd=2.7 as=0.4 ps=2.8 w=1 l=0.15
X70 a_21880_39160# a_22770_39050# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.54 as=0.168 ps=1.64 w=0.42 l=0.15
R13 uio_in[1] a_23250_39050# sky130_fd_pr__res_generic_m2 w=0.45 l=0.05
X71 a_21880_41750# a_21810_39050# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.54 as=0.168 ps=1.64 w=0.42 l=0.15
X72 a_24200_41490# a_24200_41490# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.54 as=0.168 ps=1.64 w=0.42 l=0.15
X73 ua[1] a_21880_39160# VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.55 pd=3.1 as=0.55 ps=3.1 w=1 l=0.15
X74 a_21880_41750# a_21880_41750# VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.35 pd=2.7 as=0.4 ps=2.8 w=1 l=0.15
X75 a_24200_41490# a_25610_39160# VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.35 pd=2.7 as=0.4 ps=2.8 w=1 l=0.15
X76 a_21880_39160# a_21880_39160# VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.35 pd=2.7 as=0.4 ps=2.8 w=1 l=0.15
X77 a_24200_38900# a_26090_39160# VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.35 pd=2.7 as=0.4 ps=2.8 w=1 l=0.15
X78 a_21880_39160# a_21810_39050# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.54 as=0.168 ps=1.64 w=0.42 l=0.15
X79 a_24200_38900# a_24200_38900# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.54 as=0.168 ps=1.64 w=0.42 l=0.15
R14 uio_in[7] a_21810_39050# sky130_fd_pr__res_generic_m2 w=0.45 l=0.05
R15 ui_in[1] a_25850_39160# sky130_fd_pr__res_generic_m2 w=0.45 l=0.05
C0 m2_20650_44110# uio_in[4] 0.021608f
C1 a_25370_39160# m2_27310_44110# 0.005112f
C2 a_21880_41750# VPWR 1.67321f
C3 a_24650_39160# a_25130_39160# 8.46e-19
C4 m2_28050_44110# m2_28790_44110# 0.007143f
C5 a_22530_39050# m2_20650_44110# 0.005112f
C6 a_24650_39160# a_24890_39160# 1.10933f
C7 a_21880_41750# a_25370_39160# 8.25e-21
C8 m2_19910_44110# uio_in[5] 0.021608f
C9 a_25130_39160# m2_26570_44110# 0.005112f
C10 a_21880_41750# a_25130_39160# 1.16e-20
C11 m2_27310_44110# m2_28050_44110# 0.007143f
C12 a_22290_39050# m2_19910_44110# 0.005112f
C13 a_21880_41750# a_24890_39160# 1.74e-20
C14 a_24410_39160# a_24650_39160# 1.01277f
C15 a_24890_39160# m2_25830_44110# 0.005112f
C16 a_21880_41750# a_24650_39160# 2.89e-20
C17 m2_26570_44110# m2_27310_44110# 0.007143f
C18 a_21880_41750# a_24410_39160# 0.00727f
C19 a_24650_39160# m2_25090_44110# 0.005112f
C20 m2_25830_44110# m2_26570_44110# 0.007143f
C21 a_24410_39160# m2_24350_44110# 0.005112f
C22 m2_25090_44110# m2_25830_44110# 0.007143f
C23 m2_24350_44110# m2_25090_44110# 0.007143f
C24 m2_23590_44110# m2_24350_44110# 0.006944f
C25 m2_22870_44110# m2_23590_44110# 0.007353f
C26 m2_22130_44110# m2_22870_44110# 0.007143f
C27 m2_21390_44110# m2_22130_44110# 0.007143f
C28 clk ena 0.023797f
C29 m2_20650_44110# m2_21390_44110# 0.007143f
C30 rst_n clk 0.023797f
C31 m2_19910_44110# m2_20650_44110# 0.007143f
C32 ui_in[0] rst_n 0.023797f
C33 ui_in[1] ui_in[0] 0.13387f
C34 ui_in[2] ui_in[1] 0.133768f
C35 ui_in[3] ui_in[2] 0.133458f
C36 ui_in[4] ui_in[3] 0.133435f
C37 m2_18430_44110# m2_19170_44110# 0.007143f
C38 ui_in[5] ui_in[4] 0.133252f
C39 ui_in[6] ui_in[5] 0.133228f
C40 ui_in[7] ui_in[6] 0.13321f
C41 a_21880_39160# a_24200_38900# 0.001258f
C42 a_23810_40680# a_24200_38900# 6.41e-21
C43 uio_in[0] ui_in[7] 0.132332f
C44 a_23490_39050# a_24200_38900# 0.004679f
C45 a_23810_40680# a_21880_39160# 6.87e-19
C46 VPWR ua[7] 0.010285f
C47 a_23250_39050# a_24200_38900# 1.08e-20
C48 a_23490_39050# a_21880_39160# 0.21278f
C49 uio_in[1] uio_in[0] 0.134137f
C50 a_23490_39050# uio_in[0] 0.044617f
C51 m2_19170_44110# uio_in[6] 0.021608f
C52 a_23010_39050# a_24200_38900# 6.92e-21
C53 a_23250_39050# a_21880_39160# 0.204846f
C54 a_23490_39050# a_23810_40680# 0.009378f
C55 a_26090_39160# ui_in[0] 0.049656f
C56 a_22050_39050# m2_19170_44110# 0.005112f
C57 a_22770_39050# a_24200_38900# 4.79e-21
C58 a_23010_39050# a_21880_39160# 0.204812f
C59 a_23250_39050# a_23810_40680# 8.21e-19
C60 uio_in[2] uio_in[1] 0.13321f
C61 a_26090_39160# ui_in[1] 3.52e-19
C62 a_23250_39050# uio_in[1] 0.043751f
C63 m2_18430_44110# uio_in[7] 0.021608f
C64 a_22530_39050# a_24200_38900# 4.57e-22
C65 a_22770_39050# a_21880_39160# 0.204798f
C66 a_23010_39050# a_23810_40680# 4.18e-19
C67 a_23250_39050# a_23490_39050# 1.03051f
C68 a_25850_39160# ui_in[1] 0.049419f
C69 a_26090_39160# ui_in[2] 3.3e-19
C70 a_23010_39050# uio_in[1] 0.001582f
C71 a_21810_39050# m2_18430_44110# 0.005112f
C72 a_22530_39050# a_21880_39160# 0.204791f
C73 a_22770_39050# a_23810_40680# 2.5e-19
C74 uio_in[3] uio_in[2] 0.13321f
C75 a_25850_39160# ui_in[2] 5.76e-19
C76 a_26090_39160# ui_in[3] 3.3e-19
C77 a_23010_39050# uio_in[2] 0.046102f
C78 a_21570_2680# ua[2] 0.067465f
C79 a_22290_39050# a_21880_39160# 0.204787f
C80 a_22530_39050# a_23810_40680# 1.65e-19
C81 a_23010_39050# a_23250_39050# 1.08328f
C82 m2_29530_44110# ui_in[0] 0.020029f
C83 a_25610_39160# ui_in[2] 0.051252f
C84 a_25850_39160# ui_in[3] 5.66e-19
C85 a_26090_39160# ui_in[4] 3.3e-19
C86 a_22770_39050# uio_in[2] 0.001135f
C87 a_21570_2680# ua[3] 0.297498f
C88 a_22050_39050# a_21880_39160# 0.204778f
C89 a_22290_39050# a_23810_40680# 1.17e-19
C90 uio_in[4] uio_in[3] 0.13321f
C91 a_25610_39160# ui_in[3] 6.72e-19
C92 a_25850_39160# ui_in[4] 5.53e-19
C93 a_22530_39050# uio_in[2] 8.23e-19
C94 a_22770_39050# uio_in[3] 0.047856f
C95 a_21810_39050# a_21880_39160# 0.159094f
C96 a_22770_39050# a_23010_39050# 1.19972f
C97 VPWR ui_in[4] 0.004568f
C98 m2_28790_44110# ui_in[1] 0.020255f
C99 a_25370_39160# ui_in[3] 0.049254f
C100 a_25610_39160# ui_in[4] 6.57e-19
C101 a_25850_39160# ui_in[5] 0.001163f
C102 a_22290_39050# uio_in[2] 6.38e-19
C103 a_22530_39050# uio_in[3] 8.23e-19
C104 a_24200_38900# ua[1] 0.023074f
C105 a_26090_39160# a_24200_38900# 0.143247f
C106 a_22530_39050# a_23010_39050# 1.6e-19
C107 VPWR ui_in[5] 0.004568f
C108 uio_in[5] uio_in[4] 0.13321f
C109 a_25370_39160# ui_in[4] 8.82e-19
C110 a_25610_39160# ui_in[5] 6.45e-19
C111 a_22290_39050# uio_in[3] 6.38e-19
C112 a_22530_39050# uio_in[4] 0.049358f
C113 a_21570_2680# VPWR 0.274867f
C114 a_24200_38900# ua[0] 5.38e-20
C115 a_21880_39160# ua[1] 0.072223f
C116 a_25850_39160# a_24200_38900# 0.143247f
C117 a_22290_39050# a_23010_39050# 1.13e-19
C118 a_22530_39050# a_22770_39050# 1.2778f
C119 a_24200_41490# a_23810_40680# 0.001209f
C120 VPWR ui_in[6] 0.004568f
C121 m2_28050_44110# ui_in[2] 0.02048f
C122 a_25130_39160# ui_in[4] 0.048012f
C123 a_25370_39160# ui_in[5] 8.67e-19
C124 a_22050_39050# uio_in[3] 5.15e-19
C125 a_22290_39050# uio_in[4] 6.38e-19
C126 a_24200_38900# VPWR 1.1585f
C127 a_23810_40680# ua[1] 0.273365f
C128 a_25610_39160# a_24200_38900# 0.143247f
C129 a_22290_39050# a_22770_39050# 1.23e-19
C130 a_24200_41490# a_23490_39050# 0.004011f
C131 VPWR ui_in[7] 0.004568f
C132 uio_in[6] uio_in[5] 0.13321f
C133 a_25130_39160# ui_in[5] 0.001175f
C134 a_21810_39050# uio_in[3] 2.96e-19
C135 a_22050_39050# uio_in[4] 5.15e-19
C136 a_22290_39050# uio_in[5] 0.050403f
C137 a_21880_39160# VPWR 1.5973f
C138 a_23490_39050# ua[1] 0.092903f
C139 a_23810_40680# ua[0] 0.05951f
C140 a_25370_39160# a_24200_38900# 0.143247f
C141 a_22290_39050# a_22530_39050# 1.45765f
C142 a_24200_41490# a_23250_39050# 1.08e-20
C143 a_22050_39050# a_22770_39050# 9.52e-20
C144 a_25850_39160# a_23810_40680# 9.83e-20
C145 VPWR uio_in[0] 0.004568f
C146 m2_27310_44110# ui_in[3] 0.020706f
C147 a_24890_39160# ui_in[5] 0.046777f
C148 a_25130_39160# ui_in[6] 0.004014f
C149 a_21810_39050# uio_in[4] 2.96e-19
C150 a_22050_39050# uio_in[5] 5.15e-19
C151 a_23810_40680# VPWR 0.248173f
C152 a_23250_39050# ua[1] 2.72e-19
C153 a_25130_39160# a_24200_38900# 0.143247f
C154 a_25370_39160# a_21880_39160# 4.13e-21
C155 a_24200_41490# a_23010_39050# 6.92e-21
C156 a_22050_39050# a_22530_39050# 1.18e-19
C157 a_21810_39050# a_22770_39050# 7.47e-20
C158 a_25610_39160# a_23810_40680# 1.39e-19
C159 VPWR uio_in[1] 0.004568f
C160 uio_in[7] uio_in[6] 0.13321f
C161 a_24890_39160# ui_in[6] 0.001608f
C162 a_21810_39050# uio_in[5] 2.96e-19
C163 a_22050_39050# uio_in[6] 0.051224f
C164 a_23490_39050# VPWR 0.534047f
C165 a_23010_39050# ua[1] 1.47e-19
C166 a_24890_39160# a_24200_38900# 0.143247f
C167 a_25130_39160# a_21880_39160# 5.8e-21
C168 a_24200_41490# a_22770_39050# 4.79e-21
C169 a_22050_39050# a_22290_39050# 1.64461f
C170 a_21810_39050# a_22530_39050# 9.71e-20
C171 a_25370_39160# a_23810_40680# 2.12e-19
C172 VPWR uio_in[2] 0.004568f
C173 m2_26570_44110# ui_in[4] 0.020932f
C174 a_24650_39160# ui_in[6] 0.044593f
C175 a_21810_39050# uio_in[6] 2.96e-19
C176 a_23250_39050# VPWR 0.436562f
C177 a_22770_39050# ua[1] 9.1e-20
C178 a_24650_39160# a_24200_38900# 0.143247f
C179 a_24890_39160# a_21880_39160# 8.71e-21
C180 a_24200_41490# a_22530_39050# 4.57e-22
C181 a_21810_39050# a_22290_39050# 1.06e-19
C182 a_25130_39160# a_23810_40680# 3.6e-19
C183 VPWR uio_in[3] 0.004568f
C184 a_21810_39050# uio_in[7] 0.050442f
C185 a_23010_39050# VPWR 0.439864f
C186 a_22530_39050# ua[1] 6.16e-20
C187 a_24410_39160# a_24200_38900# 0.111243f
C188 a_24650_39160# a_21880_39160# 1.44e-20
C189 a_21810_39050# a_22050_39050# 1.66539f
C190 a_24890_39160# a_23810_40680# 7.18e-19
C191 m2_25830_44110# ui_in[5] 0.021157f
C192 VPWR uio_in[4] 0.004568f
C193 a_24410_39160# ui_in[7] 0.044373f
C194 a_22770_39050# VPWR 0.445789f
C195 a_22290_39050# ua[1] 4.44e-20
C196 a_24410_39160# a_21880_39160# 0.006714f
C197 a_24650_39160# a_23810_40680# 0.001837f
C198 ua[3] ua[2] 0.038049f
C199 a_22530_39050# VPWR 0.459327f
C200 a_24410_39160# a_23810_40680# 0.049227f
C201 m2_25090_44110# ui_in[6] 0.021383f
C202 a_22290_39050# VPWR 0.478277f
C203 a_24410_39160# a_23490_39050# 0.222207f
C204 a_21880_41750# a_23810_40680# 0.002387f
C205 a_24200_41490# ua[1] 0.019982f
C206 a_22050_39050# VPWR 0.510229f
C207 a_26090_39160# a_24200_41490# 0.215989f
C208 a_21880_41750# a_23490_39050# 0.229552f
C209 VPWR ua[2] 0.206244f
C210 m2_24350_44110# ui_in[7] 0.021608f
C211 a_26090_39160# ua[1] 1.8e-19
C212 a_24200_41490# ua[0] 0.001164f
C213 a_21810_39050# VPWR 0.87516f
C214 a_25850_39160# a_24200_41490# 0.221092f
C215 a_21880_41750# a_23250_39050# 0.221622f
C216 VPWR ua[3] 0.346539f
C217 a_25850_39160# ua[1] 1.8e-19
C218 a_26090_39160# ua[0] 0.100513f
C219 a_24200_41490# VPWR 1.2358f
C220 a_25610_39160# a_24200_41490# 0.21981f
C221 a_25850_39160# a_26090_39160# 1.68469f
C222 a_21880_41750# a_23010_39050# 0.221772f
C223 m2_23590_44110# uio_in[0] 0.021608f
C224 VPWR ua[1] 0.709125f
C225 a_25610_39160# ua[1] 1.8e-19
C226 a_25850_39160# ua[0] 0.05653f
C227 m2_19170_44110# m2_19910_44110# 0.007143f
C228 a_26090_39160# VPWR 0.90977f
C229 a_25370_39160# a_24200_41490# 0.220682f
C230 a_25610_39160# a_26090_39160# 1.54e-19
C231 a_21880_41750# a_22770_39050# 0.222103f
C232 VPWR ua[0] 0.765277f
C233 a_23490_39050# m2_23590_44110# 0.005112f
C234 a_25370_39160# ua[1] 1.8e-19
C235 a_25610_39160# ua[0] 0.055424f
C236 a_25850_39160# VPWR 0.567946f
C237 a_25130_39160# a_24200_41490# 0.219289f
C238 a_25370_39160# a_26090_39160# 1.28e-19
C239 a_25610_39160# a_25850_39160# 1.89777f
C240 a_21880_41750# a_22530_39050# 0.222316f
C241 m2_22870_44110# uio_in[1] 0.021608f
C242 a_25130_39160# ua[1] 1.8e-19
C243 a_25370_39160# ua[0] 0.055026f
C244 a_25610_39160# VPWR 0.553411f
C245 a_26090_39160# m2_29530_44110# 0.005112f
C246 a_24890_39160# a_24200_41490# 0.220228f
C247 a_25130_39160# a_26090_39160# 1.13e-19
C248 a_25370_39160# a_25850_39160# 1.49e-19
C249 a_21880_41750# a_22290_39050# 0.2225f
C250 a_23250_39050# m2_22870_44110# 0.005112f
C251 a_24890_39160# ua[1] 1.8e-19
C252 a_25130_39160# ua[0] 0.055076f
C253 a_25370_39160# VPWR 0.537607f
C254 a_24650_39160# a_24200_41490# 0.219087f
C255 a_25130_39160# a_25850_39160# 1.34e-19
C256 a_25370_39160# a_25610_39160# 1.3709f
C257 a_21880_41750# a_22050_39050# 0.222751f
C258 m2_22130_44110# uio_in[2] 0.021608f
C259 a_25850_39160# m2_28790_44110# 0.005112f
C260 a_24650_39160# ua[1] 1.8e-19
C261 a_24890_39160# ua[0] 0.055733f
C262 a_25130_39160# VPWR 0.527069f
C263 a_24410_39160# a_24200_41490# 0.18266f
C264 a_24890_39160# a_25850_39160# 3.05e-19
C265 a_25130_39160# a_25610_39160# 1.56e-19
C266 a_21880_41750# a_21810_39050# 0.16944f
C267 a_23010_39050# m2_22130_44110# 0.005112f
C268 a_24650_39160# ua[0] 0.06855f
C269 a_24410_39160# ua[1] 0.093209f
C270 a_24890_39160# VPWR 0.520247f
C271 a_24890_39160# a_25610_39160# 1.23e-19
C272 a_25130_39160# a_25370_39160# 1.31698f
C273 a_21880_41750# a_24200_41490# 0.001258f
C274 m2_21390_44110# uio_in[3] 0.021608f
C275 a_25610_39160# m2_28050_44110# 0.005112f
C276 a_24410_39160# ua[0] 0.111655f
C277 a_21880_41750# ua[1] 0.071522f
C278 a_24650_39160# VPWR 0.531904f
C279 a_24890_39160# a_25370_39160# 1.78e-19
C280 m2_28790_44110# m2_29530_44110# 0.007143f
C281 a_22770_39050# m2_21390_44110# 0.005112f
C282 a_24410_39160# VPWR 0.663104f
C283 a_24890_39160# a_25130_39160# 1.21119f
C284 ua[4] VGND 0.122428f
C285 ua[5] VGND 0.122428f
C286 ua[6] VGND 0.122428f
C287 ua[7] VGND 0.111009f
C288 ena VGND 0.073297f
C289 clk VGND 0.0487f
C290 rst_n VGND 0.0487f
C291 ui_in[0] VGND 0.350951f
C292 ui_in[1] VGND 0.234234f
C293 ui_in[2] VGND 0.230502f
C294 ui_in[3] VGND 0.230704f
C295 ui_in[4] VGND 0.223397f
C296 ui_in[5] VGND 0.22191f
C297 ui_in[6] VGND 0.220814f
C298 ui_in[7] VGND 0.223871f
C299 uio_in[0] VGND 0.225466f
C300 uio_in[1] VGND 0.224179f
C301 uio_in[2] VGND 0.221286f
C302 uio_in[3] VGND 0.219592f
C303 uio_in[4] VGND 0.218871f
C304 uio_in[5] VGND 0.224716f
C305 uio_in[6] VGND 0.224366f
C306 uio_in[7] VGND 0.362103f
C307 ua[2] VGND 1.67217f
C308 ua[3] VGND 3.44482f
C309 ua[1] VGND 18.018312f
C310 ua[0] VGND 18.881802f
C311 VPWR VGND 78.8463f
C312 m2_29530_44110# VGND 0.049454f $ **FLOATING
C313 m2_28790_44110# VGND 0.040694f $ **FLOATING
C314 m2_28050_44110# VGND 0.040694f $ **FLOATING
C315 m2_27310_44110# VGND 0.040694f $ **FLOATING
C316 m2_26570_44110# VGND 0.040694f $ **FLOATING
C317 m2_25830_44110# VGND 0.040694f $ **FLOATING
C318 m2_25090_44110# VGND 0.040694f $ **FLOATING
C319 m2_24350_44110# VGND 0.040877f $ **FLOATING
C320 m2_23590_44110# VGND 0.040687f $ **FLOATING
C321 m2_22870_44110# VGND 0.040504f $ **FLOATING
C322 m2_22130_44110# VGND 0.040694f $ **FLOATING
C323 m2_21390_44110# VGND 0.040694f $ **FLOATING
C324 m2_20650_44110# VGND 0.040694f $ **FLOATING
C325 m2_19910_44110# VGND 0.040694f $ **FLOATING
C326 m2_19170_44110# VGND 0.040694f $ **FLOATING
C327 m2_18430_44110# VGND 0.049454f $ **FLOATING
C328 a_21570_2680# VGND 0.711945f
C329 a_24200_38900# VGND 2.73692f
C330 a_21880_39160# VGND 1.994f
C331 a_23810_40680# VGND 0.712389f
C332 a_23490_39050# VGND 1.66046f
C333 a_23250_39050# VGND 1.41306f
C334 a_23010_39050# VGND 1.54891f
C335 a_22770_39050# VGND 1.64741f
C336 a_22530_39050# VGND 1.73515f
C337 a_22290_39050# VGND 1.80588f
C338 a_22050_39050# VGND 1.90533f
C339 a_21810_39050# VGND 3.17095f
C340 a_24200_41490# VGND 2.66092f
C341 a_26090_39160# VGND 2.90456f
C342 a_25850_39160# VGND 1.70481f
C343 a_25610_39160# VGND 1.62106f
C344 a_25370_39160# VGND 1.57552f
C345 a_25130_39160# VGND 1.47461f
C346 a_24890_39160# VGND 1.37037f
C347 a_24650_39160# VGND 1.22953f
C348 a_24410_39160# VGND 1.37675f
C349 a_21880_41750# VGND 1.92325f


.ends

* set gnd and power
Vgnd VGND 0 0
Vdd VPWR VGND 1.8

* create pulse
* Vin A VGND pulse(0 1.8 1p 10p 10p 1n 2n)
* Isource A VGND pulse(-0.001 0.001 0 500p 500p 500p 2n)

* Vin0 X0 VGND pulse(0 1.8 1p 10p 10p 1n 2n)
* Vin1 X1 VGND 0
* Vin2 Y0 VGND pulse(0 1.8 500p 10p 10p 1n 2n)
* Vin3 Y1 VGND 0
* .tran 10e-12 2e-09 0e-00

*   112233
*  5050505
* 01210121
* 000011112222

* pulse(0 1.8  5n 10p 10p 10n 20n)
* pulse(0 1.8 10n 10p 10p 10n 20n)
* pulse(0 1.8 20n 10p 10p 20n 40n)
* pulse(0 1.8  1p 10p 10p 20n 40n)

VinY0 Y0 VGND pulse(1.8 0  20n 10p 10p 100n 160n)
VinY1 Y1 VGND pulse(1.8 0  40n 10p 10p 100n 160n)
VinY2 Y2 VGND pulse(1.8 0  60n 10p 10p 100n 160n)
VinY3 Y3 VGND pulse(1.8 0  80n 10p 10p 100n 160n)
VinY4 Y4 VGND pulse(1.8 0 100n 10p 10p 100n 160n)
VinY5 Y5 VGND 1.8
VinY6 Y6 VGND 1.8
VinY7 Y7 VGND 1.8

VinX0 X0 VGND pulse(0 1.8  5n 10p 10p 20n 40n)
VinX1 X1 VGND pulse(0 1.8 10n 10p 10p 20n 40n)
VinX2 X2 VGND pulse(0 1.8 15n 10p 10p 20n 40n)
VinX3 X3 VGND pulse(0 1.8 20n 10p 10p 20n 40n)
VinX4 X4 VGND 0
VinX5 X5 VGND 0
VinX6 X6 VGND 0
VinX7 X7 VGND 0

.tran 10e-12 12e-08 0e-00

.control
run
set color0 = white
set color1 = black
plot X0 X1 X2 X3
plot Y0 Y1 Y2 Y3 Y4
plot Out
plot i(Vdd)
.endc
