magic
tech sky130A
magscale 1 2
timestamp 1713286768
<< nwell >>
rect 11240 42960 11600 43350
<< nmos >>
rect 11400 42720 11430 42804
<< pmos >>
rect 11400 43000 11430 43200
<< ndiff >>
rect 11320 42780 11400 42804
rect 11320 42740 11340 42780
rect 11380 42740 11400 42780
rect 11320 42720 11400 42740
rect 11430 42780 11520 42804
rect 11430 42740 11450 42780
rect 11490 42740 11520 42780
rect 11430 42720 11520 42740
<< pdiff >>
rect 11320 43170 11400 43200
rect 11320 43030 11340 43170
rect 11380 43030 11400 43170
rect 11320 43000 11400 43030
rect 11430 43170 11520 43200
rect 11430 43030 11450 43170
rect 11490 43030 11520 43170
rect 11430 43000 11520 43030
<< ndiffc >>
rect 11340 42740 11380 42780
rect 11450 42740 11490 42780
<< pdiffc >>
rect 11340 43030 11380 43170
rect 11450 43030 11490 43170
<< psubdiff >>
rect 11300 42610 11330 42650
rect 11370 42610 11400 42650
rect 11460 42610 11490 42650
rect 11530 42610 11560 42650
<< nsubdiff >>
rect 11300 43270 11330 43310
rect 11370 43270 11400 43310
rect 11460 43270 11490 43310
rect 11530 43270 11560 43310
<< psubdiffcont >>
rect 11330 42610 11370 42650
rect 11490 42610 11530 42650
<< nsubdiffcont >>
rect 11330 43270 11370 43310
rect 11490 43270 11530 43310
<< poly >>
rect 11400 43200 11430 43240
rect 11400 42930 11430 43000
rect 11320 42910 11430 42930
rect 11320 42870 11340 42910
rect 11380 42870 11430 42910
rect 11320 42850 11430 42870
rect 11400 42804 11430 42850
rect 11400 42680 11430 42720
<< polycont >>
rect 11340 42870 11380 42910
<< locali >>
rect 11000 43310 11550 43330
rect 11000 43270 11020 43310
rect 11060 43270 11330 43310
rect 11370 43270 11490 43310
rect 11530 43270 11550 43310
rect 11000 43250 11550 43270
rect 11320 43170 11380 43250
rect 11320 43030 11340 43170
rect 11320 43000 11380 43030
rect 11450 43170 11510 43200
rect 11490 43030 11510 43170
rect 11450 42910 11510 43030
rect 11250 42870 11340 42910
rect 11380 42870 11400 42910
rect 11450 42870 11550 42910
rect 11320 42780 11380 42800
rect 11320 42740 11340 42780
rect 11320 42670 11380 42740
rect 11450 42780 11510 42870
rect 11490 42740 11510 42780
rect 11450 42720 11510 42740
rect 11010 42650 11550 42670
rect 11010 42610 11030 42650
rect 11070 42610 11330 42650
rect 11370 42610 11490 42650
rect 11530 42610 11550 42650
rect 11010 42590 11550 42610
<< viali >>
rect 11020 43270 11060 43310
rect 11030 42610 11070 42650
<< metal1 >>
rect 10740 43380 11140 43390
rect 10740 43200 10750 43380
rect 10930 43310 11140 43380
rect 10930 43270 11020 43310
rect 11060 43270 11140 43310
rect 10930 43200 11140 43270
rect 10740 43190 11140 43200
rect 10740 42710 11140 42720
rect 10740 42530 10750 42710
rect 10930 42650 11140 42710
rect 10930 42610 11030 42650
rect 11070 42610 11140 42650
rect 10930 42530 11140 42610
rect 10740 42520 11140 42530
<< via1 >>
rect 10750 43200 10930 43380
rect 10750 42530 10930 42710
<< metal2 >>
rect 10540 43380 10940 43390
rect 10540 43200 10550 43380
rect 10730 43200 10750 43380
rect 10930 43200 10940 43380
rect 10540 43190 10940 43200
rect 10540 42710 10940 42720
rect 10540 42530 10550 42710
rect 10730 42530 10750 42710
rect 10930 42530 10940 42710
rect 10540 42520 10940 42530
<< via2 >>
rect 10550 43200 10730 43380
rect 10550 42530 10730 42710
<< metal3 >>
rect 8898 43460 10740 43470
rect 8898 43180 8910 43460
rect 9190 43380 10740 43460
rect 9190 43200 10550 43380
rect 10730 43200 10740 43380
rect 9190 43180 10740 43200
rect 8898 43170 10740 43180
rect 10340 42710 10740 42720
rect 10340 42530 10350 42710
rect 10530 42530 10550 42710
rect 10730 42530 10740 42710
rect 10340 42520 10740 42530
rect 201 22427 8861 22725
<< via3 >>
rect 8910 43180 9190 43460
rect 10350 42530 10530 42710
<< metal4 >>
rect 798 44952 858 45152
rect 1534 44952 1594 45152
rect 2270 44952 2330 45152
rect 3006 44952 3066 45152
rect 3742 44952 3802 45152
rect 4478 44952 4538 45152
rect 5214 44952 5274 45152
rect 5950 44952 6010 45152
rect 6686 44952 6746 45152
rect 7422 44952 7482 45152
rect 8158 44952 8218 45152
rect 8894 44952 8954 45152
rect 9630 44952 9690 45152
rect 10366 44952 10426 45152
rect 11102 44952 11162 45152
rect 11838 44952 11898 45152
rect 12574 44952 12634 45152
rect 13310 44952 13370 45152
rect 14046 44952 14106 45152
rect 14782 44952 14842 45152
rect 15518 44952 15578 45152
rect 16254 44952 16314 45152
rect 16990 44952 17050 45152
rect 17726 44952 17786 45152
rect 18462 44952 18522 45152
rect 19198 44952 19258 45152
rect 19934 44952 19994 45152
rect 20670 44952 20730 45152
rect 21406 44952 21466 45152
rect 22142 44952 22202 45152
rect 22878 44952 22938 45152
rect 23614 44952 23674 45152
rect 24350 44952 24410 45152
rect 25086 44952 25146 45152
rect 25822 44952 25882 45152
rect 26558 44952 26618 45152
rect 27294 44952 27354 45152
rect 28030 44952 28090 45152
rect 28766 44952 28826 45152
rect 29502 44952 29562 45152
rect 30238 44952 30298 45152
rect 30974 44952 31034 45152
rect 31710 44952 31770 45152
rect 200 43470 500 44152
rect 200 43460 9198 43470
rect 200 43180 8910 43460
rect 9190 43180 9198 43460
rect 200 43170 9198 43180
rect 200 1000 500 43170
rect 9800 42798 10100 44152
rect 9800 42710 10540 42798
rect 9800 42530 10350 42710
rect 10530 42530 10540 42710
rect 9800 42498 10540 42530
rect 9800 1000 10100 42498
rect 400 0 520 200
rect 4816 0 4936 200
rect 9232 0 9352 200
rect 13648 0 13768 200
rect 18064 0 18184 200
rect 22480 0 22600 200
rect 26896 0 27016 200
rect 31312 0 31432 200
<< labels >>
flabel metal4 s 30974 44952 31034 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 31710 44952 31770 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 30238 44952 30298 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 31312 0 31432 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26896 0 27016 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22480 0 22600 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18064 0 18184 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 13648 0 13768 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 9232 0 9352 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 4816 0 4936 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 400 0 520 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 29502 44952 29562 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 28030 44952 28090 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 27294 44952 27354 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 25822 44952 25882 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 25086 44952 25146 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23614 44952 23674 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22878 44952 22938 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21406 44952 21466 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 20670 44952 20730 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19198 44952 19258 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 18462 44952 18522 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 5950 44952 6010 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 5214 44952 5274 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 4478 44952 4538 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 3742 44952 3802 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 3006 44952 3066 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 2270 44952 2330 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 1534 44952 1594 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 798 44952 858 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 11838 44952 11898 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 10366 44952 10426 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 9630 44952 9690 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 8158 44952 8218 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 7422 44952 7482 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 16990 44952 17050 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 16254 44952 16314 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 14782 44952 14842 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 14046 44952 14106 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 12574 44952 12634 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 200 1000 500 44152 1 FreeSans 2 0 0 0 VPWR
port 51 nsew power bidirectional
flabel metal4 9800 1000 10100 44152 1 FreeSans 2 0 0 0 VGND
port 52 nsew ground bidirectional
rlabel locali 11250 42870 11290 42910 1 A
rlabel locali 11510 42870 11550 42910 1 Y
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
