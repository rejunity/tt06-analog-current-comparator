magic
tech sky130A
magscale 1 2
timestamp 1713389596
<< nwell >>
rect 12870 42970 13600 43350
<< nmos >>
rect 13070 42710 13100 42794
rect 13400 42710 13430 42794
<< pmos >>
rect 13070 43010 13100 43210
rect 13400 43010 13430 43210
<< ndiff >>
rect 12980 42770 13070 42794
rect 12980 42730 13010 42770
rect 13050 42730 13070 42770
rect 12980 42710 13070 42730
rect 13100 42770 13180 42794
rect 13100 42730 13120 42770
rect 13160 42730 13180 42770
rect 13100 42710 13180 42730
rect 13320 42770 13400 42794
rect 13320 42730 13340 42770
rect 13380 42730 13400 42770
rect 13320 42710 13400 42730
rect 13430 42770 13520 42794
rect 13430 42730 13450 42770
rect 13490 42730 13520 42770
rect 13430 42710 13520 42730
<< pdiff >>
rect 12910 43180 13070 43210
rect 12910 43040 12930 43180
rect 12970 43040 13070 43180
rect 12910 43010 13070 43040
rect 13100 43180 13180 43210
rect 13100 43040 13120 43180
rect 13160 43040 13180 43180
rect 13100 43010 13180 43040
rect 13320 43180 13400 43210
rect 13320 43040 13340 43180
rect 13380 43040 13400 43180
rect 13320 43010 13400 43040
rect 13430 43180 13520 43210
rect 13430 43040 13450 43180
rect 13490 43040 13520 43180
rect 13430 43010 13520 43040
<< ndiffc >>
rect 13010 42730 13050 42770
rect 13120 42730 13160 42770
rect 13340 42730 13380 42770
rect 13450 42730 13490 42770
<< pdiffc >>
rect 12930 43040 12970 43180
rect 13120 43040 13160 43180
rect 13340 43040 13380 43180
rect 13450 43040 13490 43180
<< psubdiff >>
rect 12980 42610 13010 42650
rect 13050 42610 13080 42650
rect 13140 42610 13170 42650
rect 13210 42610 13240 42650
rect 13300 42610 13330 42650
rect 13370 42610 13400 42650
rect 13460 42610 13490 42650
rect 13530 42610 13560 42650
<< nsubdiff >>
rect 12980 43270 13010 43310
rect 13050 43270 13080 43310
rect 13140 43270 13170 43310
rect 13210 43270 13240 43310
rect 13300 43270 13330 43310
rect 13370 43270 13400 43310
rect 13460 43270 13490 43310
rect 13530 43270 13560 43310
<< psubdiffcont >>
rect 13010 42610 13050 42650
rect 13170 42610 13210 42650
rect 13330 42610 13370 42650
rect 13490 42610 13530 42650
<< nsubdiffcont >>
rect 13010 43270 13050 43310
rect 13170 43270 13210 43310
rect 13330 43270 13370 43310
rect 13490 43270 13530 43310
<< poly >>
rect 13070 43210 13100 43240
rect 13400 43210 13430 43240
rect 13070 42890 13100 43010
rect 13400 42970 13430 43010
rect 13320 42960 13430 42970
rect 13320 42920 13340 42960
rect 13380 42920 13430 42960
rect 13320 42910 13430 42920
rect 13070 42880 13280 42890
rect 13070 42840 13220 42880
rect 13260 42840 13280 42880
rect 13070 42830 13280 42840
rect 13070 42794 13100 42830
rect 13400 42794 13430 42910
rect 13070 42680 13100 42710
rect 13400 42680 13430 42710
<< polycont >>
rect 13340 42920 13380 42960
rect 13220 42840 13260 42880
<< locali >>
rect 11000 43310 13550 43330
rect 11000 43270 11020 43310
rect 11060 43270 13010 43310
rect 13050 43270 13170 43310
rect 13210 43270 13330 43310
rect 13370 43270 13490 43310
rect 13530 43270 13550 43310
rect 11000 43250 13550 43270
rect 12930 43180 12970 43210
rect 12930 42670 12970 43040
rect 13010 42770 13050 43250
rect 13010 42710 13050 42730
rect 13120 43180 13160 43210
rect 13120 42960 13160 43040
rect 13320 43180 13380 43250
rect 13320 43040 13340 43180
rect 13320 43010 13380 43040
rect 13450 43180 13510 43210
rect 13490 43040 13510 43180
rect 13120 42920 13340 42960
rect 13380 42920 13400 42960
rect 13450 42920 13510 43040
rect 13120 42770 13160 42920
rect 13450 42880 13550 42920
rect 13200 42840 13220 42880
rect 13260 42840 13510 42880
rect 13120 42710 13160 42730
rect 13320 42770 13380 42790
rect 13320 42730 13340 42770
rect 13320 42670 13380 42730
rect 13450 42770 13510 42840
rect 13490 42730 13510 42770
rect 13450 42710 13510 42730
rect 11010 42650 13550 42670
rect 11010 42610 11030 42650
rect 11070 42610 13010 42650
rect 13050 42610 13170 42650
rect 13210 42610 13330 42650
rect 13370 42610 13490 42650
rect 13530 42610 13550 42650
rect 11010 42590 13550 42610
<< viali >>
rect 11020 43270 11060 43310
rect 11030 42610 11070 42650
<< metal1 >>
rect 10740 43380 11140 43390
rect 10740 43200 10750 43380
rect 10930 43310 11140 43380
rect 10930 43270 11020 43310
rect 11060 43270 11140 43310
rect 10930 43200 11140 43270
rect 10740 43190 11140 43200
rect 10740 42710 11140 42720
rect 10740 42530 10750 42710
rect 10930 42650 11140 42710
rect 10930 42610 11030 42650
rect 11070 42610 11140 42650
rect 10930 42530 11140 42610
rect 10740 42520 11140 42530
<< via1 >>
rect 10750 43200 10930 43380
rect 10750 42530 10930 42710
<< metal2 >>
rect 10540 43380 10940 43390
rect 10540 43200 10550 43380
rect 10730 43200 10750 43380
rect 10930 43200 10940 43380
rect 10540 43190 10940 43200
rect 10540 42710 10940 42720
rect 10540 42530 10550 42710
rect 10730 42530 10750 42710
rect 10930 42530 10940 42710
rect 10540 42520 10940 42530
<< via2 >>
rect 10550 43200 10730 43380
rect 10550 42530 10730 42710
<< metal3 >>
rect 8898 43460 10740 43470
rect 8898 43180 8910 43460
rect 9190 43380 10740 43460
rect 9190 43200 10550 43380
rect 10730 43200 10740 43380
rect 9190 43180 10740 43200
rect 8898 43170 10740 43180
rect 10340 42710 10740 42720
rect 10340 42530 10350 42710
rect 10530 42530 10550 42710
rect 10730 42530 10740 42710
rect 10340 42520 10740 42530
rect 201 22427 8861 22725
<< via3 >>
rect 8910 43180 9190 43460
rect 10350 42530 10530 42710
<< metal4 >>
rect 798 44952 858 45152
rect 1534 44952 1594 45152
rect 2270 44952 2330 45152
rect 3006 44952 3066 45152
rect 3742 44952 3802 45152
rect 4478 44952 4538 45152
rect 5214 44952 5274 45152
rect 5950 44952 6010 45152
rect 6686 44952 6746 45152
rect 7422 44952 7482 45152
rect 8158 44952 8218 45152
rect 8894 44952 8954 45152
rect 9630 44952 9690 45152
rect 10366 44952 10426 45152
rect 11102 44952 11162 45152
rect 11838 44952 11898 45152
rect 12574 44952 12634 45152
rect 13310 44952 13370 45152
rect 14046 44952 14106 45152
rect 14782 44952 14842 45152
rect 15518 44952 15578 45152
rect 16254 44952 16314 45152
rect 16990 44952 17050 45152
rect 17726 44952 17786 45152
rect 18462 44952 18522 45152
rect 19198 44952 19258 45152
rect 19934 44952 19994 45152
rect 20670 44952 20730 45152
rect 21406 44952 21466 45152
rect 22142 44952 22202 45152
rect 22878 44952 22938 45152
rect 23614 44952 23674 45152
rect 24350 44952 24410 45152
rect 25086 44952 25146 45152
rect 25822 44952 25882 45152
rect 26558 44952 26618 45152
rect 27294 44952 27354 45152
rect 28030 44952 28090 45152
rect 28766 44952 28826 45152
rect 29502 44952 29562 45152
rect 30238 44952 30298 45152
rect 30974 44952 31034 45152
rect 31710 44952 31770 45152
rect 200 43470 500 44152
rect 200 43460 9198 43470
rect 200 43180 8910 43460
rect 9190 43180 9198 43460
rect 200 43170 9198 43180
rect 200 1000 500 43170
rect 9800 42798 10100 44152
rect 9800 42710 10540 42798
rect 9800 42530 10350 42710
rect 10530 42530 10540 42710
rect 9800 42498 10540 42530
rect 9800 1000 10100 42498
rect 400 0 520 200
rect 4816 0 4936 200
rect 9232 0 9352 200
rect 13648 0 13768 200
rect 18064 0 18184 200
rect 22480 0 22600 200
rect 26896 0 27016 200
rect 31312 0 31432 200
<< labels >>
flabel metal4 s 30974 44952 31034 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 31710 44952 31770 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 30238 44952 30298 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 31312 0 31432 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26896 0 27016 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22480 0 22600 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18064 0 18184 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 13648 0 13768 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 9232 0 9352 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 4816 0 4936 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 400 0 520 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 29502 44952 29562 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 28030 44952 28090 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 27294 44952 27354 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 25822 44952 25882 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 25086 44952 25146 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23614 44952 23674 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22878 44952 22938 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21406 44952 21466 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 20670 44952 20730 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19198 44952 19258 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 18462 44952 18522 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 5950 44952 6010 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 5214 44952 5274 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 4478 44952 4538 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 3742 44952 3802 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 3006 44952 3066 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 2270 44952 2330 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 1534 44952 1594 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 798 44952 858 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 10366 44952 10426 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 9630 44952 9690 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 8158 44952 8218 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 7422 44952 7482 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 16990 44952 17050 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 16254 44952 16314 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 14782 44952 14842 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 14046 44952 14106 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 12574 44952 12634 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 11838 44952 11898 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 200 1000 500 44152 1 FreeSans 2 0 0 0 VPWR
port 51 nsew power bidirectional
flabel metal4 9800 1000 10100 44152 1 FreeSans 2 0 0 0 VGND
port 52 nsew ground bidirectional
rlabel locali 13510 42880 13550 42920 1 Y
rlabel locali 13250 42920 13290 42960 1 A
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
