magic
tech sky130A
magscale 1 2
timestamp 1713482736
<< nwell >>
rect 21660 41810 26360 42190
rect 23610 40970 24660 41350
rect 12870 38970 13600 39350
rect 21660 39220 26360 39600
<< nmos >>
rect 21880 41520 21910 41604
rect 22120 41520 22150 41604
rect 22360 41520 22390 41604
rect 22600 41520 22630 41604
rect 22840 41520 22870 41604
rect 23080 41520 23110 41604
rect 23320 41520 23350 41604
rect 23560 41520 23590 41604
rect 24200 41520 24230 41604
rect 24480 41520 24510 41604
rect 24720 41520 24750 41604
rect 24960 41520 24990 41604
rect 25200 41520 25230 41604
rect 25440 41520 25470 41604
rect 25680 41520 25710 41604
rect 25920 41520 25950 41604
rect 26160 41520 26190 41604
rect 23810 40710 23840 40794
rect 24140 40710 24170 40794
rect 24400 40710 24430 40794
rect 21880 38930 21910 39014
rect 22120 38930 22150 39014
rect 22360 38930 22390 39014
rect 22600 38930 22630 39014
rect 22840 38930 22870 39014
rect 23080 38930 23110 39014
rect 23320 38930 23350 39014
rect 23560 38930 23590 39014
rect 24200 38930 24230 39014
rect 24480 38930 24510 39014
rect 24720 38930 24750 39014
rect 24960 38930 24990 39014
rect 25200 38930 25230 39014
rect 25440 38930 25470 39014
rect 25680 38930 25710 39014
rect 25920 38930 25950 39014
rect 26160 38930 26190 39014
rect 13070 38710 13100 38794
rect 13400 38710 13430 38794
<< pmos >>
rect 21880 41850 21910 42050
rect 22120 41850 22150 42050
rect 22360 41850 22390 42050
rect 22600 41850 22630 42050
rect 22840 41850 22870 42050
rect 23080 41850 23110 42050
rect 23320 41850 23350 42050
rect 23560 41850 23590 42050
rect 23880 41850 23910 42050
rect 24480 41850 24510 42050
rect 24720 41850 24750 42050
rect 24960 41850 24990 42050
rect 25200 41850 25230 42050
rect 25440 41850 25470 42050
rect 25680 41850 25710 42050
rect 25920 41850 25950 42050
rect 26160 41850 26190 42050
rect 23810 41010 23840 41210
rect 24140 41010 24170 41210
rect 24400 41010 24430 41210
rect 21880 39260 21910 39460
rect 22120 39260 22150 39460
rect 22360 39260 22390 39460
rect 22600 39260 22630 39460
rect 22840 39260 22870 39460
rect 23080 39260 23110 39460
rect 23320 39260 23350 39460
rect 23560 39260 23590 39460
rect 23880 39260 23910 39460
rect 24480 39260 24510 39460
rect 24720 39260 24750 39460
rect 24960 39260 24990 39460
rect 25200 39260 25230 39460
rect 25440 39260 25470 39460
rect 25680 39260 25710 39460
rect 25920 39260 25950 39460
rect 26160 39260 26190 39460
rect 13070 39010 13100 39210
rect 13400 39010 13430 39210
<< ndiff >>
rect 21800 41580 21880 41604
rect 21800 41540 21820 41580
rect 21860 41540 21880 41580
rect 21800 41520 21880 41540
rect 21910 41580 21980 41604
rect 21910 41540 21930 41580
rect 21970 41540 21980 41580
rect 21910 41520 21980 41540
rect 22040 41580 22120 41604
rect 22040 41540 22060 41580
rect 22100 41540 22120 41580
rect 22040 41520 22120 41540
rect 22150 41580 22220 41604
rect 22150 41540 22170 41580
rect 22210 41540 22220 41580
rect 22150 41520 22220 41540
rect 22280 41580 22360 41604
rect 22280 41540 22300 41580
rect 22340 41540 22360 41580
rect 22280 41520 22360 41540
rect 22390 41580 22460 41604
rect 22390 41540 22410 41580
rect 22450 41540 22460 41580
rect 22390 41520 22460 41540
rect 22520 41580 22600 41604
rect 22520 41540 22540 41580
rect 22580 41540 22600 41580
rect 22520 41520 22600 41540
rect 22630 41580 22700 41604
rect 22630 41540 22650 41580
rect 22690 41540 22700 41580
rect 22630 41520 22700 41540
rect 22760 41580 22840 41604
rect 22760 41540 22780 41580
rect 22820 41540 22840 41580
rect 22760 41520 22840 41540
rect 22870 41580 22940 41604
rect 22870 41540 22890 41580
rect 22930 41540 22940 41580
rect 22870 41520 22940 41540
rect 23000 41580 23080 41604
rect 23000 41540 23020 41580
rect 23060 41540 23080 41580
rect 23000 41520 23080 41540
rect 23110 41580 23180 41604
rect 23110 41540 23130 41580
rect 23170 41540 23180 41580
rect 23110 41520 23180 41540
rect 23240 41580 23320 41604
rect 23240 41540 23260 41580
rect 23300 41540 23320 41580
rect 23240 41520 23320 41540
rect 23350 41580 23420 41604
rect 23350 41540 23370 41580
rect 23410 41540 23420 41580
rect 23350 41520 23420 41540
rect 23480 41580 23560 41604
rect 23480 41540 23500 41580
rect 23540 41540 23560 41580
rect 23480 41520 23560 41540
rect 23590 41580 23660 41604
rect 23590 41540 23610 41580
rect 23650 41540 23660 41580
rect 23590 41520 23660 41540
rect 24090 41580 24200 41604
rect 24090 41540 24100 41580
rect 24180 41540 24200 41580
rect 24090 41520 24200 41540
rect 24230 41580 24340 41604
rect 24230 41540 24250 41580
rect 24330 41540 24340 41580
rect 24230 41520 24340 41540
rect 24400 41580 24480 41604
rect 24400 41540 24420 41580
rect 24460 41540 24480 41580
rect 24400 41520 24480 41540
rect 24510 41580 24580 41604
rect 24510 41540 24530 41580
rect 24570 41540 24580 41580
rect 24510 41520 24580 41540
rect 24640 41580 24720 41604
rect 24640 41540 24660 41580
rect 24700 41540 24720 41580
rect 24640 41520 24720 41540
rect 24750 41580 24820 41604
rect 24750 41540 24770 41580
rect 24810 41540 24820 41580
rect 24750 41520 24820 41540
rect 24880 41580 24960 41604
rect 24880 41540 24900 41580
rect 24940 41540 24960 41580
rect 24880 41520 24960 41540
rect 24990 41580 25060 41604
rect 24990 41540 25010 41580
rect 25050 41540 25060 41580
rect 24990 41520 25060 41540
rect 25120 41580 25200 41604
rect 25120 41540 25140 41580
rect 25180 41540 25200 41580
rect 25120 41520 25200 41540
rect 25230 41580 25300 41604
rect 25230 41540 25250 41580
rect 25290 41540 25300 41580
rect 25230 41520 25300 41540
rect 25360 41580 25440 41604
rect 25360 41540 25380 41580
rect 25420 41540 25440 41580
rect 25360 41520 25440 41540
rect 25470 41580 25540 41604
rect 25470 41540 25490 41580
rect 25530 41540 25540 41580
rect 25470 41520 25540 41540
rect 25600 41580 25680 41604
rect 25600 41540 25620 41580
rect 25660 41540 25680 41580
rect 25600 41520 25680 41540
rect 25710 41580 25780 41604
rect 25710 41540 25730 41580
rect 25770 41540 25780 41580
rect 25710 41520 25780 41540
rect 25840 41580 25920 41604
rect 25840 41540 25860 41580
rect 25900 41540 25920 41580
rect 25840 41520 25920 41540
rect 25950 41580 26020 41604
rect 25950 41540 25970 41580
rect 26010 41540 26020 41580
rect 25950 41520 26020 41540
rect 26080 41580 26160 41604
rect 26080 41540 26100 41580
rect 26140 41540 26160 41580
rect 26080 41520 26160 41540
rect 26190 41580 26260 41604
rect 26190 41540 26210 41580
rect 26250 41540 26260 41580
rect 26190 41520 26260 41540
rect 23720 40770 23810 40794
rect 23720 40730 23750 40770
rect 23790 40730 23810 40770
rect 23720 40710 23810 40730
rect 23840 40770 23920 40794
rect 23840 40730 23860 40770
rect 23900 40730 23920 40770
rect 23840 40710 23920 40730
rect 24060 40770 24140 40794
rect 24060 40730 24080 40770
rect 24120 40730 24140 40770
rect 24060 40710 24140 40730
rect 24170 40770 24260 40794
rect 24170 40730 24190 40770
rect 24230 40730 24260 40770
rect 24170 40710 24260 40730
rect 24320 40770 24400 40794
rect 24320 40730 24340 40770
rect 24380 40730 24400 40770
rect 24320 40710 24400 40730
rect 24430 40770 24520 40794
rect 24430 40730 24450 40770
rect 24490 40730 24520 40770
rect 24430 40710 24520 40730
rect 21800 38990 21880 39014
rect 21800 38950 21820 38990
rect 21860 38950 21880 38990
rect 21800 38930 21880 38950
rect 21910 38990 21980 39014
rect 21910 38950 21930 38990
rect 21970 38950 21980 38990
rect 21910 38930 21980 38950
rect 22040 38990 22120 39014
rect 22040 38950 22060 38990
rect 22100 38950 22120 38990
rect 22040 38930 22120 38950
rect 22150 38990 22220 39014
rect 22150 38950 22170 38990
rect 22210 38950 22220 38990
rect 22150 38930 22220 38950
rect 22280 38990 22360 39014
rect 22280 38950 22300 38990
rect 22340 38950 22360 38990
rect 22280 38930 22360 38950
rect 22390 38990 22460 39014
rect 22390 38950 22410 38990
rect 22450 38950 22460 38990
rect 22390 38930 22460 38950
rect 22520 38990 22600 39014
rect 22520 38950 22540 38990
rect 22580 38950 22600 38990
rect 22520 38930 22600 38950
rect 22630 38990 22700 39014
rect 22630 38950 22650 38990
rect 22690 38950 22700 38990
rect 22630 38930 22700 38950
rect 22760 38990 22840 39014
rect 22760 38950 22780 38990
rect 22820 38950 22840 38990
rect 22760 38930 22840 38950
rect 22870 38990 22940 39014
rect 22870 38950 22890 38990
rect 22930 38950 22940 38990
rect 22870 38930 22940 38950
rect 23000 38990 23080 39014
rect 23000 38950 23020 38990
rect 23060 38950 23080 38990
rect 23000 38930 23080 38950
rect 23110 38990 23180 39014
rect 23110 38950 23130 38990
rect 23170 38950 23180 38990
rect 23110 38930 23180 38950
rect 23240 38990 23320 39014
rect 23240 38950 23260 38990
rect 23300 38950 23320 38990
rect 23240 38930 23320 38950
rect 23350 38990 23420 39014
rect 23350 38950 23370 38990
rect 23410 38950 23420 38990
rect 23350 38930 23420 38950
rect 23480 38990 23560 39014
rect 23480 38950 23500 38990
rect 23540 38950 23560 38990
rect 23480 38930 23560 38950
rect 23590 38990 23660 39014
rect 23590 38950 23610 38990
rect 23650 38950 23660 38990
rect 23590 38930 23660 38950
rect 24090 38990 24200 39014
rect 24090 38950 24100 38990
rect 24180 38950 24200 38990
rect 24090 38930 24200 38950
rect 24230 38990 24340 39014
rect 24230 38950 24250 38990
rect 24330 38950 24340 38990
rect 24230 38930 24340 38950
rect 24400 38990 24480 39014
rect 24400 38950 24420 38990
rect 24460 38950 24480 38990
rect 24400 38930 24480 38950
rect 24510 38990 24580 39014
rect 24510 38950 24530 38990
rect 24570 38950 24580 38990
rect 24510 38930 24580 38950
rect 24640 38990 24720 39014
rect 24640 38950 24660 38990
rect 24700 38950 24720 38990
rect 24640 38930 24720 38950
rect 24750 38990 24820 39014
rect 24750 38950 24770 38990
rect 24810 38950 24820 38990
rect 24750 38930 24820 38950
rect 24880 38990 24960 39014
rect 24880 38950 24900 38990
rect 24940 38950 24960 38990
rect 24880 38930 24960 38950
rect 24990 38990 25060 39014
rect 24990 38950 25010 38990
rect 25050 38950 25060 38990
rect 24990 38930 25060 38950
rect 25120 38990 25200 39014
rect 25120 38950 25140 38990
rect 25180 38950 25200 38990
rect 25120 38930 25200 38950
rect 25230 38990 25300 39014
rect 25230 38950 25250 38990
rect 25290 38950 25300 38990
rect 25230 38930 25300 38950
rect 25360 38990 25440 39014
rect 25360 38950 25380 38990
rect 25420 38950 25440 38990
rect 25360 38930 25440 38950
rect 25470 38990 25540 39014
rect 25470 38950 25490 38990
rect 25530 38950 25540 38990
rect 25470 38930 25540 38950
rect 25600 38990 25680 39014
rect 25600 38950 25620 38990
rect 25660 38950 25680 38990
rect 25600 38930 25680 38950
rect 25710 38990 25780 39014
rect 25710 38950 25730 38990
rect 25770 38950 25780 38990
rect 25710 38930 25780 38950
rect 25840 38990 25920 39014
rect 25840 38950 25860 38990
rect 25900 38950 25920 38990
rect 25840 38930 25920 38950
rect 25950 38990 26020 39014
rect 25950 38950 25970 38990
rect 26010 38950 26020 38990
rect 25950 38930 26020 38950
rect 26080 38990 26160 39014
rect 26080 38950 26100 38990
rect 26140 38950 26160 38990
rect 26080 38930 26160 38950
rect 26190 38990 26260 39014
rect 26190 38950 26210 38990
rect 26250 38950 26260 38990
rect 26190 38930 26260 38950
rect 12980 38770 13070 38794
rect 12980 38730 13010 38770
rect 13050 38730 13070 38770
rect 12980 38710 13070 38730
rect 13100 38770 13180 38794
rect 13100 38730 13120 38770
rect 13160 38730 13180 38770
rect 13100 38710 13180 38730
rect 13320 38770 13400 38794
rect 13320 38730 13340 38770
rect 13380 38730 13400 38770
rect 13320 38710 13400 38730
rect 13430 38770 13520 38794
rect 13430 38730 13450 38770
rect 13490 38730 13520 38770
rect 13430 38710 13520 38730
<< pdiff >>
rect 21800 42020 21880 42050
rect 21800 41880 21820 42020
rect 21860 41880 21880 42020
rect 21800 41850 21880 41880
rect 21910 42020 21980 42050
rect 21910 41880 21930 42020
rect 21970 41880 21980 42020
rect 21910 41850 21980 41880
rect 22040 42020 22120 42050
rect 22040 41880 22060 42020
rect 22100 41880 22120 42020
rect 22040 41850 22120 41880
rect 22150 42020 22220 42050
rect 22150 41880 22170 42020
rect 22210 41880 22220 42020
rect 22150 41850 22220 41880
rect 22280 42020 22360 42050
rect 22280 41880 22300 42020
rect 22340 41880 22360 42020
rect 22280 41850 22360 41880
rect 22390 42020 22460 42050
rect 22390 41880 22410 42020
rect 22450 41880 22460 42020
rect 22390 41850 22460 41880
rect 22520 42020 22600 42050
rect 22520 41880 22540 42020
rect 22580 41880 22600 42020
rect 22520 41850 22600 41880
rect 22630 42020 22700 42050
rect 22630 41880 22650 42020
rect 22690 41880 22700 42020
rect 22630 41850 22700 41880
rect 22760 42020 22840 42050
rect 22760 41880 22780 42020
rect 22820 41880 22840 42020
rect 22760 41850 22840 41880
rect 22870 42020 22940 42050
rect 22870 41880 22890 42020
rect 22930 41880 22940 42020
rect 22870 41850 22940 41880
rect 23000 42020 23080 42050
rect 23000 41880 23020 42020
rect 23060 41880 23080 42020
rect 23000 41850 23080 41880
rect 23110 42020 23180 42050
rect 23110 41880 23130 42020
rect 23170 41880 23180 42020
rect 23110 41850 23180 41880
rect 23240 42020 23320 42050
rect 23240 41880 23260 42020
rect 23300 41880 23320 42020
rect 23240 41850 23320 41880
rect 23350 42020 23420 42050
rect 23350 41880 23370 42020
rect 23410 41880 23420 42020
rect 23350 41850 23420 41880
rect 23480 42020 23560 42050
rect 23480 41880 23500 42020
rect 23540 41880 23560 42020
rect 23480 41850 23560 41880
rect 23590 42020 23660 42050
rect 23590 41880 23610 42020
rect 23650 41880 23660 42020
rect 23590 41850 23660 41880
rect 23770 42020 23880 42050
rect 23770 41880 23780 42020
rect 23860 41880 23880 42020
rect 23770 41850 23880 41880
rect 23910 42020 24020 42050
rect 23910 41880 23930 42020
rect 24010 41880 24020 42020
rect 23910 41850 24020 41880
rect 24400 42020 24480 42050
rect 24400 41880 24420 42020
rect 24460 41880 24480 42020
rect 24400 41850 24480 41880
rect 24510 42020 24580 42050
rect 24510 41880 24530 42020
rect 24570 41880 24580 42020
rect 24510 41850 24580 41880
rect 24640 42020 24720 42050
rect 24640 41880 24660 42020
rect 24700 41880 24720 42020
rect 24640 41850 24720 41880
rect 24750 42020 24820 42050
rect 24750 41880 24770 42020
rect 24810 41880 24820 42020
rect 24750 41850 24820 41880
rect 24880 42020 24960 42050
rect 24880 41880 24900 42020
rect 24940 41880 24960 42020
rect 24880 41850 24960 41880
rect 24990 42020 25060 42050
rect 24990 41880 25010 42020
rect 25050 41880 25060 42020
rect 24990 41850 25060 41880
rect 25120 42020 25200 42050
rect 25120 41880 25140 42020
rect 25180 41880 25200 42020
rect 25120 41850 25200 41880
rect 25230 42020 25300 42050
rect 25230 41880 25250 42020
rect 25290 41880 25300 42020
rect 25230 41850 25300 41880
rect 25360 42020 25440 42050
rect 25360 41880 25380 42020
rect 25420 41880 25440 42020
rect 25360 41850 25440 41880
rect 25470 42020 25540 42050
rect 25470 41880 25490 42020
rect 25530 41880 25540 42020
rect 25470 41850 25540 41880
rect 25600 42020 25680 42050
rect 25600 41880 25620 42020
rect 25660 41880 25680 42020
rect 25600 41850 25680 41880
rect 25710 42020 25780 42050
rect 25710 41880 25730 42020
rect 25770 41880 25780 42020
rect 25710 41850 25780 41880
rect 25840 42020 25920 42050
rect 25840 41880 25860 42020
rect 25900 41880 25920 42020
rect 25840 41850 25920 41880
rect 25950 42020 26020 42050
rect 25950 41880 25970 42020
rect 26010 41880 26020 42020
rect 25950 41850 26020 41880
rect 26080 42020 26160 42050
rect 26080 41880 26100 42020
rect 26140 41880 26160 42020
rect 26080 41850 26160 41880
rect 26190 42020 26260 42050
rect 26190 41880 26210 42020
rect 26250 41880 26260 42020
rect 26190 41850 26260 41880
rect 23650 41180 23810 41210
rect 23650 41040 23670 41180
rect 23710 41040 23810 41180
rect 23650 41010 23810 41040
rect 23840 41180 23920 41210
rect 23840 41040 23860 41180
rect 23900 41040 23920 41180
rect 23840 41010 23920 41040
rect 24060 41180 24140 41210
rect 24060 41040 24080 41180
rect 24120 41040 24140 41180
rect 24060 41010 24140 41040
rect 24170 41180 24260 41210
rect 24170 41040 24190 41180
rect 24230 41040 24260 41180
rect 24170 41010 24260 41040
rect 24320 41180 24400 41210
rect 24320 41040 24340 41180
rect 24380 41040 24400 41180
rect 24320 41010 24400 41040
rect 24430 41180 24520 41210
rect 24430 41040 24450 41180
rect 24490 41040 24520 41180
rect 24430 41010 24520 41040
rect 21800 39430 21880 39460
rect 21800 39290 21820 39430
rect 21860 39290 21880 39430
rect 21800 39260 21880 39290
rect 21910 39430 21980 39460
rect 21910 39290 21930 39430
rect 21970 39290 21980 39430
rect 21910 39260 21980 39290
rect 22040 39430 22120 39460
rect 22040 39290 22060 39430
rect 22100 39290 22120 39430
rect 22040 39260 22120 39290
rect 22150 39430 22220 39460
rect 22150 39290 22170 39430
rect 22210 39290 22220 39430
rect 22150 39260 22220 39290
rect 22280 39430 22360 39460
rect 22280 39290 22300 39430
rect 22340 39290 22360 39430
rect 22280 39260 22360 39290
rect 22390 39430 22460 39460
rect 22390 39290 22410 39430
rect 22450 39290 22460 39430
rect 22390 39260 22460 39290
rect 22520 39430 22600 39460
rect 22520 39290 22540 39430
rect 22580 39290 22600 39430
rect 22520 39260 22600 39290
rect 22630 39430 22700 39460
rect 22630 39290 22650 39430
rect 22690 39290 22700 39430
rect 22630 39260 22700 39290
rect 22760 39430 22840 39460
rect 22760 39290 22780 39430
rect 22820 39290 22840 39430
rect 22760 39260 22840 39290
rect 22870 39430 22940 39460
rect 22870 39290 22890 39430
rect 22930 39290 22940 39430
rect 22870 39260 22940 39290
rect 23000 39430 23080 39460
rect 23000 39290 23020 39430
rect 23060 39290 23080 39430
rect 23000 39260 23080 39290
rect 23110 39430 23180 39460
rect 23110 39290 23130 39430
rect 23170 39290 23180 39430
rect 23110 39260 23180 39290
rect 23240 39430 23320 39460
rect 23240 39290 23260 39430
rect 23300 39290 23320 39430
rect 23240 39260 23320 39290
rect 23350 39430 23420 39460
rect 23350 39290 23370 39430
rect 23410 39290 23420 39430
rect 23350 39260 23420 39290
rect 23480 39430 23560 39460
rect 23480 39290 23500 39430
rect 23540 39290 23560 39430
rect 23480 39260 23560 39290
rect 23590 39430 23660 39460
rect 23590 39290 23610 39430
rect 23650 39290 23660 39430
rect 23590 39260 23660 39290
rect 23770 39430 23880 39460
rect 23770 39290 23780 39430
rect 23860 39290 23880 39430
rect 23770 39260 23880 39290
rect 23910 39430 24020 39460
rect 23910 39290 23930 39430
rect 24010 39290 24020 39430
rect 23910 39260 24020 39290
rect 24400 39430 24480 39460
rect 24400 39290 24420 39430
rect 24460 39290 24480 39430
rect 24400 39260 24480 39290
rect 24510 39430 24580 39460
rect 24510 39290 24530 39430
rect 24570 39290 24580 39430
rect 24510 39260 24580 39290
rect 24640 39430 24720 39460
rect 24640 39290 24660 39430
rect 24700 39290 24720 39430
rect 24640 39260 24720 39290
rect 24750 39430 24820 39460
rect 24750 39290 24770 39430
rect 24810 39290 24820 39430
rect 24750 39260 24820 39290
rect 24880 39430 24960 39460
rect 24880 39290 24900 39430
rect 24940 39290 24960 39430
rect 24880 39260 24960 39290
rect 24990 39430 25060 39460
rect 24990 39290 25010 39430
rect 25050 39290 25060 39430
rect 24990 39260 25060 39290
rect 25120 39430 25200 39460
rect 25120 39290 25140 39430
rect 25180 39290 25200 39430
rect 25120 39260 25200 39290
rect 25230 39430 25300 39460
rect 25230 39290 25250 39430
rect 25290 39290 25300 39430
rect 25230 39260 25300 39290
rect 25360 39430 25440 39460
rect 25360 39290 25380 39430
rect 25420 39290 25440 39430
rect 25360 39260 25440 39290
rect 25470 39430 25540 39460
rect 25470 39290 25490 39430
rect 25530 39290 25540 39430
rect 25470 39260 25540 39290
rect 25600 39430 25680 39460
rect 25600 39290 25620 39430
rect 25660 39290 25680 39430
rect 25600 39260 25680 39290
rect 25710 39430 25780 39460
rect 25710 39290 25730 39430
rect 25770 39290 25780 39430
rect 25710 39260 25780 39290
rect 25840 39430 25920 39460
rect 25840 39290 25860 39430
rect 25900 39290 25920 39430
rect 25840 39260 25920 39290
rect 25950 39430 26020 39460
rect 25950 39290 25970 39430
rect 26010 39290 26020 39430
rect 25950 39260 26020 39290
rect 26080 39430 26160 39460
rect 26080 39290 26100 39430
rect 26140 39290 26160 39430
rect 26080 39260 26160 39290
rect 26190 39430 26260 39460
rect 26190 39290 26210 39430
rect 26250 39290 26260 39430
rect 26190 39260 26260 39290
rect 12910 39180 13070 39210
rect 12910 39040 12930 39180
rect 12970 39040 13070 39180
rect 12910 39010 13070 39040
rect 13100 39180 13180 39210
rect 13100 39040 13120 39180
rect 13160 39040 13180 39180
rect 13100 39010 13180 39040
rect 13320 39180 13400 39210
rect 13320 39040 13340 39180
rect 13380 39040 13400 39180
rect 13320 39010 13400 39040
rect 13430 39180 13520 39210
rect 13430 39040 13450 39180
rect 13490 39040 13520 39180
rect 13430 39010 13520 39040
<< ndiffc >>
rect 21820 41540 21860 41580
rect 21930 41540 21970 41580
rect 22060 41540 22100 41580
rect 22170 41540 22210 41580
rect 22300 41540 22340 41580
rect 22410 41540 22450 41580
rect 22540 41540 22580 41580
rect 22650 41540 22690 41580
rect 22780 41540 22820 41580
rect 22890 41540 22930 41580
rect 23020 41540 23060 41580
rect 23130 41540 23170 41580
rect 23260 41540 23300 41580
rect 23370 41540 23410 41580
rect 23500 41540 23540 41580
rect 23610 41540 23650 41580
rect 24100 41540 24180 41580
rect 24250 41540 24330 41580
rect 24420 41540 24460 41580
rect 24530 41540 24570 41580
rect 24660 41540 24700 41580
rect 24770 41540 24810 41580
rect 24900 41540 24940 41580
rect 25010 41540 25050 41580
rect 25140 41540 25180 41580
rect 25250 41540 25290 41580
rect 25380 41540 25420 41580
rect 25490 41540 25530 41580
rect 25620 41540 25660 41580
rect 25730 41540 25770 41580
rect 25860 41540 25900 41580
rect 25970 41540 26010 41580
rect 26100 41540 26140 41580
rect 26210 41540 26250 41580
rect 23750 40730 23790 40770
rect 23860 40730 23900 40770
rect 24080 40730 24120 40770
rect 24190 40730 24230 40770
rect 24340 40730 24380 40770
rect 24450 40730 24490 40770
rect 21820 38950 21860 38990
rect 21930 38950 21970 38990
rect 22060 38950 22100 38990
rect 22170 38950 22210 38990
rect 22300 38950 22340 38990
rect 22410 38950 22450 38990
rect 22540 38950 22580 38990
rect 22650 38950 22690 38990
rect 22780 38950 22820 38990
rect 22890 38950 22930 38990
rect 23020 38950 23060 38990
rect 23130 38950 23170 38990
rect 23260 38950 23300 38990
rect 23370 38950 23410 38990
rect 23500 38950 23540 38990
rect 23610 38950 23650 38990
rect 24100 38950 24180 38990
rect 24250 38950 24330 38990
rect 24420 38950 24460 38990
rect 24530 38950 24570 38990
rect 24660 38950 24700 38990
rect 24770 38950 24810 38990
rect 24900 38950 24940 38990
rect 25010 38950 25050 38990
rect 25140 38950 25180 38990
rect 25250 38950 25290 38990
rect 25380 38950 25420 38990
rect 25490 38950 25530 38990
rect 25620 38950 25660 38990
rect 25730 38950 25770 38990
rect 25860 38950 25900 38990
rect 25970 38950 26010 38990
rect 26100 38950 26140 38990
rect 26210 38950 26250 38990
rect 13010 38730 13050 38770
rect 13120 38730 13160 38770
rect 13340 38730 13380 38770
rect 13450 38730 13490 38770
<< pdiffc >>
rect 21820 41880 21860 42020
rect 21930 41880 21970 42020
rect 22060 41880 22100 42020
rect 22170 41880 22210 42020
rect 22300 41880 22340 42020
rect 22410 41880 22450 42020
rect 22540 41880 22580 42020
rect 22650 41880 22690 42020
rect 22780 41880 22820 42020
rect 22890 41880 22930 42020
rect 23020 41880 23060 42020
rect 23130 41880 23170 42020
rect 23260 41880 23300 42020
rect 23370 41880 23410 42020
rect 23500 41880 23540 42020
rect 23610 41880 23650 42020
rect 23780 41880 23860 42020
rect 23930 41880 24010 42020
rect 24420 41880 24460 42020
rect 24530 41880 24570 42020
rect 24660 41880 24700 42020
rect 24770 41880 24810 42020
rect 24900 41880 24940 42020
rect 25010 41880 25050 42020
rect 25140 41880 25180 42020
rect 25250 41880 25290 42020
rect 25380 41880 25420 42020
rect 25490 41880 25530 42020
rect 25620 41880 25660 42020
rect 25730 41880 25770 42020
rect 25860 41880 25900 42020
rect 25970 41880 26010 42020
rect 26100 41880 26140 42020
rect 26210 41880 26250 42020
rect 23670 41040 23710 41180
rect 23860 41040 23900 41180
rect 24080 41040 24120 41180
rect 24190 41040 24230 41180
rect 24340 41040 24380 41180
rect 24450 41040 24490 41180
rect 21820 39290 21860 39430
rect 21930 39290 21970 39430
rect 22060 39290 22100 39430
rect 22170 39290 22210 39430
rect 22300 39290 22340 39430
rect 22410 39290 22450 39430
rect 22540 39290 22580 39430
rect 22650 39290 22690 39430
rect 22780 39290 22820 39430
rect 22890 39290 22930 39430
rect 23020 39290 23060 39430
rect 23130 39290 23170 39430
rect 23260 39290 23300 39430
rect 23370 39290 23410 39430
rect 23500 39290 23540 39430
rect 23610 39290 23650 39430
rect 23780 39290 23860 39430
rect 23930 39290 24010 39430
rect 24420 39290 24460 39430
rect 24530 39290 24570 39430
rect 24660 39290 24700 39430
rect 24770 39290 24810 39430
rect 24900 39290 24940 39430
rect 25010 39290 25050 39430
rect 25140 39290 25180 39430
rect 25250 39290 25290 39430
rect 25380 39290 25420 39430
rect 25490 39290 25530 39430
rect 25620 39290 25660 39430
rect 25730 39290 25770 39430
rect 25860 39290 25900 39430
rect 25970 39290 26010 39430
rect 26100 39290 26140 39430
rect 26210 39290 26250 39430
rect 12930 39040 12970 39180
rect 13120 39040 13160 39180
rect 13340 39040 13380 39180
rect 13450 39040 13490 39180
<< psubdiff >>
rect 21700 41420 21730 41460
rect 21770 41420 21800 41460
rect 21860 41420 21890 41460
rect 21930 41420 21960 41460
rect 22020 41420 22050 41460
rect 22090 41420 22120 41460
rect 22180 41420 22210 41460
rect 22250 41420 22280 41460
rect 22340 41420 22370 41460
rect 22410 41420 22440 41460
rect 22500 41420 22530 41460
rect 22570 41420 22600 41460
rect 22660 41420 22690 41460
rect 22730 41420 22760 41460
rect 22820 41420 22850 41460
rect 22890 41420 22920 41460
rect 22980 41420 23010 41460
rect 23050 41420 23080 41460
rect 23140 41420 23170 41460
rect 23210 41420 23240 41460
rect 23300 41420 23330 41460
rect 23370 41420 23400 41460
rect 23460 41420 23490 41460
rect 23530 41420 23560 41460
rect 23620 41420 23650 41460
rect 23690 41420 23720 41460
rect 24140 41420 24170 41460
rect 24210 41420 24240 41460
rect 24300 41420 24330 41460
rect 24370 41420 24400 41460
rect 24460 41420 24490 41460
rect 24530 41420 24560 41460
rect 24620 41420 24650 41460
rect 24690 41420 24720 41460
rect 24780 41420 24810 41460
rect 24850 41420 24880 41460
rect 24940 41420 24970 41460
rect 25010 41420 25040 41460
rect 25100 41420 25130 41460
rect 25170 41420 25200 41460
rect 25260 41420 25290 41460
rect 25330 41420 25360 41460
rect 25420 41420 25450 41460
rect 25490 41420 25520 41460
rect 25580 41420 25610 41460
rect 25650 41420 25680 41460
rect 25740 41420 25770 41460
rect 25810 41420 25840 41460
rect 25900 41420 25930 41460
rect 25970 41420 26000 41460
rect 26060 41420 26090 41460
rect 26130 41420 26160 41460
rect 26220 41420 26250 41460
rect 26290 41420 26320 41460
rect 23720 40610 23750 40650
rect 23790 40610 23820 40650
rect 23880 40610 23910 40650
rect 23950 40610 23980 40650
rect 24040 40610 24070 40650
rect 24110 40610 24140 40650
rect 24200 40610 24230 40650
rect 24270 40610 24300 40650
rect 24360 40610 24390 40650
rect 24430 40610 24460 40650
rect 24520 40610 24550 40650
rect 24590 40610 24620 40650
rect 21700 38830 21730 38870
rect 21770 38830 21800 38870
rect 21860 38830 21890 38870
rect 21930 38830 21960 38870
rect 22020 38830 22050 38870
rect 22090 38830 22120 38870
rect 22180 38830 22210 38870
rect 22250 38830 22280 38870
rect 22340 38830 22370 38870
rect 22410 38830 22440 38870
rect 22500 38830 22530 38870
rect 22570 38830 22600 38870
rect 22660 38830 22690 38870
rect 22730 38830 22760 38870
rect 22820 38830 22850 38870
rect 22890 38830 22920 38870
rect 22980 38830 23010 38870
rect 23050 38830 23080 38870
rect 23140 38830 23170 38870
rect 23210 38830 23240 38870
rect 23300 38830 23330 38870
rect 23370 38830 23400 38870
rect 23460 38830 23490 38870
rect 23530 38830 23560 38870
rect 23620 38830 23650 38870
rect 23690 38830 23720 38870
rect 24140 38830 24170 38870
rect 24210 38830 24240 38870
rect 24300 38830 24330 38870
rect 24370 38830 24400 38870
rect 24460 38830 24490 38870
rect 24530 38830 24560 38870
rect 24620 38830 24650 38870
rect 24690 38830 24720 38870
rect 24780 38830 24810 38870
rect 24850 38830 24880 38870
rect 24940 38830 24970 38870
rect 25010 38830 25040 38870
rect 25100 38830 25130 38870
rect 25170 38830 25200 38870
rect 25260 38830 25290 38870
rect 25330 38830 25360 38870
rect 25420 38830 25450 38870
rect 25490 38830 25520 38870
rect 25580 38830 25610 38870
rect 25650 38830 25680 38870
rect 25740 38830 25770 38870
rect 25810 38830 25840 38870
rect 25900 38830 25930 38870
rect 25970 38830 26000 38870
rect 26060 38830 26090 38870
rect 26130 38830 26160 38870
rect 26220 38830 26250 38870
rect 26290 38830 26320 38870
rect 12980 38610 13010 38650
rect 13050 38610 13080 38650
rect 13140 38610 13170 38650
rect 13210 38610 13240 38650
rect 13300 38610 13330 38650
rect 13370 38610 13400 38650
rect 13460 38610 13490 38650
rect 13530 38610 13560 38650
<< nsubdiff >>
rect 21700 42110 21730 42150
rect 21770 42110 21800 42150
rect 21860 42110 21890 42150
rect 21930 42110 21960 42150
rect 22020 42110 22050 42150
rect 22090 42110 22120 42150
rect 22180 42110 22210 42150
rect 22250 42110 22280 42150
rect 22340 42110 22370 42150
rect 22410 42110 22440 42150
rect 22500 42110 22530 42150
rect 22570 42110 22600 42150
rect 22660 42110 22690 42150
rect 22730 42110 22760 42150
rect 22820 42110 22850 42150
rect 22890 42110 22920 42150
rect 22980 42110 23010 42150
rect 23050 42110 23080 42150
rect 23140 42110 23170 42150
rect 23210 42110 23240 42150
rect 23300 42110 23330 42150
rect 23370 42110 23400 42150
rect 23460 42110 23490 42150
rect 23530 42110 23560 42150
rect 23620 42110 23650 42150
rect 23690 42110 23720 42150
rect 23780 42110 23810 42150
rect 23850 42110 23880 42150
rect 23940 42110 23970 42150
rect 24010 42110 24040 42150
rect 24300 42110 24330 42150
rect 24370 42110 24400 42150
rect 24460 42110 24490 42150
rect 24530 42110 24560 42150
rect 24620 42110 24650 42150
rect 24690 42110 24720 42150
rect 24780 42110 24810 42150
rect 24850 42110 24880 42150
rect 24940 42110 24970 42150
rect 25010 42110 25040 42150
rect 25100 42110 25130 42150
rect 25170 42110 25200 42150
rect 25260 42110 25290 42150
rect 25330 42110 25360 42150
rect 25420 42110 25450 42150
rect 25490 42110 25520 42150
rect 25580 42110 25610 42150
rect 25650 42110 25680 42150
rect 25740 42110 25770 42150
rect 25810 42110 25840 42150
rect 25900 42110 25930 42150
rect 25970 42110 26000 42150
rect 26060 42110 26090 42150
rect 26130 42110 26160 42150
rect 26220 42110 26250 42150
rect 26290 42110 26320 42150
rect 23720 41270 23750 41310
rect 23790 41270 23820 41310
rect 23880 41270 23910 41310
rect 23950 41270 23980 41310
rect 24040 41270 24070 41310
rect 24110 41270 24140 41310
rect 24200 41270 24230 41310
rect 24270 41270 24300 41310
rect 24360 41270 24390 41310
rect 24430 41270 24460 41310
rect 24520 41270 24550 41310
rect 24590 41270 24620 41310
rect 21700 39520 21730 39560
rect 21770 39520 21800 39560
rect 21860 39520 21890 39560
rect 21930 39520 21960 39560
rect 22020 39520 22050 39560
rect 22090 39520 22120 39560
rect 22180 39520 22210 39560
rect 22250 39520 22280 39560
rect 22340 39520 22370 39560
rect 22410 39520 22440 39560
rect 22500 39520 22530 39560
rect 22570 39520 22600 39560
rect 22660 39520 22690 39560
rect 22730 39520 22760 39560
rect 22820 39520 22850 39560
rect 22890 39520 22920 39560
rect 22980 39520 23010 39560
rect 23050 39520 23080 39560
rect 23140 39520 23170 39560
rect 23210 39520 23240 39560
rect 23300 39520 23330 39560
rect 23370 39520 23400 39560
rect 23460 39520 23490 39560
rect 23530 39520 23560 39560
rect 23620 39520 23650 39560
rect 23690 39520 23720 39560
rect 23780 39520 23810 39560
rect 23850 39520 23880 39560
rect 23940 39520 23970 39560
rect 24010 39520 24040 39560
rect 24300 39520 24330 39560
rect 24370 39520 24400 39560
rect 24460 39520 24490 39560
rect 24530 39520 24560 39560
rect 24620 39520 24650 39560
rect 24690 39520 24720 39560
rect 24780 39520 24810 39560
rect 24850 39520 24880 39560
rect 24940 39520 24970 39560
rect 25010 39520 25040 39560
rect 25100 39520 25130 39560
rect 25170 39520 25200 39560
rect 25260 39520 25290 39560
rect 25330 39520 25360 39560
rect 25420 39520 25450 39560
rect 25490 39520 25520 39560
rect 25580 39520 25610 39560
rect 25650 39520 25680 39560
rect 25740 39520 25770 39560
rect 25810 39520 25840 39560
rect 25900 39520 25930 39560
rect 25970 39520 26000 39560
rect 26060 39520 26090 39560
rect 26130 39520 26160 39560
rect 26220 39520 26250 39560
rect 26290 39520 26320 39560
rect 12980 39270 13010 39310
rect 13050 39270 13080 39310
rect 13140 39270 13170 39310
rect 13210 39270 13240 39310
rect 13300 39270 13330 39310
rect 13370 39270 13400 39310
rect 13460 39270 13490 39310
rect 13530 39270 13560 39310
<< psubdiffcont >>
rect 21730 41420 21770 41460
rect 21890 41420 21930 41460
rect 22050 41420 22090 41460
rect 22210 41420 22250 41460
rect 22370 41420 22410 41460
rect 22530 41420 22570 41460
rect 22690 41420 22730 41460
rect 22850 41420 22890 41460
rect 23010 41420 23050 41460
rect 23170 41420 23210 41460
rect 23330 41420 23370 41460
rect 23490 41420 23530 41460
rect 23650 41420 23690 41460
rect 24170 41420 24210 41460
rect 24330 41420 24370 41460
rect 24490 41420 24530 41460
rect 24650 41420 24690 41460
rect 24810 41420 24850 41460
rect 24970 41420 25010 41460
rect 25130 41420 25170 41460
rect 25290 41420 25330 41460
rect 25450 41420 25490 41460
rect 25610 41420 25650 41460
rect 25770 41420 25810 41460
rect 25930 41420 25970 41460
rect 26090 41420 26130 41460
rect 26250 41420 26290 41460
rect 23750 40610 23790 40650
rect 23910 40610 23950 40650
rect 24070 40610 24110 40650
rect 24230 40610 24270 40650
rect 24390 40610 24430 40650
rect 24550 40610 24590 40650
rect 21730 38830 21770 38870
rect 21890 38830 21930 38870
rect 22050 38830 22090 38870
rect 22210 38830 22250 38870
rect 22370 38830 22410 38870
rect 22530 38830 22570 38870
rect 22690 38830 22730 38870
rect 22850 38830 22890 38870
rect 23010 38830 23050 38870
rect 23170 38830 23210 38870
rect 23330 38830 23370 38870
rect 23490 38830 23530 38870
rect 23650 38830 23690 38870
rect 24170 38830 24210 38870
rect 24330 38830 24370 38870
rect 24490 38830 24530 38870
rect 24650 38830 24690 38870
rect 24810 38830 24850 38870
rect 24970 38830 25010 38870
rect 25130 38830 25170 38870
rect 25290 38830 25330 38870
rect 25450 38830 25490 38870
rect 25610 38830 25650 38870
rect 25770 38830 25810 38870
rect 25930 38830 25970 38870
rect 26090 38830 26130 38870
rect 26250 38830 26290 38870
rect 13010 38610 13050 38650
rect 13170 38610 13210 38650
rect 13330 38610 13370 38650
rect 13490 38610 13530 38650
<< nsubdiffcont >>
rect 21730 42110 21770 42150
rect 21890 42110 21930 42150
rect 22050 42110 22090 42150
rect 22210 42110 22250 42150
rect 22370 42110 22410 42150
rect 22530 42110 22570 42150
rect 22690 42110 22730 42150
rect 22850 42110 22890 42150
rect 23010 42110 23050 42150
rect 23170 42110 23210 42150
rect 23330 42110 23370 42150
rect 23490 42110 23530 42150
rect 23650 42110 23690 42150
rect 23810 42110 23850 42150
rect 23970 42110 24010 42150
rect 24330 42110 24370 42150
rect 24490 42110 24530 42150
rect 24650 42110 24690 42150
rect 24810 42110 24850 42150
rect 24970 42110 25010 42150
rect 25130 42110 25170 42150
rect 25290 42110 25330 42150
rect 25450 42110 25490 42150
rect 25610 42110 25650 42150
rect 25770 42110 25810 42150
rect 25930 42110 25970 42150
rect 26090 42110 26130 42150
rect 26250 42110 26290 42150
rect 23750 41270 23790 41310
rect 23910 41270 23950 41310
rect 24070 41270 24110 41310
rect 24230 41270 24270 41310
rect 24390 41270 24430 41310
rect 24550 41270 24590 41310
rect 21730 39520 21770 39560
rect 21890 39520 21930 39560
rect 22050 39520 22090 39560
rect 22210 39520 22250 39560
rect 22370 39520 22410 39560
rect 22530 39520 22570 39560
rect 22690 39520 22730 39560
rect 22850 39520 22890 39560
rect 23010 39520 23050 39560
rect 23170 39520 23210 39560
rect 23330 39520 23370 39560
rect 23490 39520 23530 39560
rect 23650 39520 23690 39560
rect 23810 39520 23850 39560
rect 23970 39520 24010 39560
rect 24330 39520 24370 39560
rect 24490 39520 24530 39560
rect 24650 39520 24690 39560
rect 24810 39520 24850 39560
rect 24970 39520 25010 39560
rect 25130 39520 25170 39560
rect 25290 39520 25330 39560
rect 25450 39520 25490 39560
rect 25610 39520 25650 39560
rect 25770 39520 25810 39560
rect 25930 39520 25970 39560
rect 26090 39520 26130 39560
rect 26250 39520 26290 39560
rect 13010 39270 13050 39310
rect 13170 39270 13210 39310
rect 13330 39270 13370 39310
rect 13490 39270 13530 39310
<< poly >>
rect 21880 42050 21910 42080
rect 22120 42050 22150 42080
rect 22360 42050 22390 42080
rect 22600 42050 22630 42080
rect 22840 42050 22870 42080
rect 23080 42050 23110 42080
rect 23320 42050 23350 42080
rect 23560 42050 23590 42080
rect 23880 42050 23910 42080
rect 24480 42050 24510 42080
rect 24720 42050 24750 42080
rect 24960 42050 24990 42080
rect 25200 42050 25230 42080
rect 25440 42050 25470 42080
rect 25680 42050 25710 42080
rect 25920 42050 25950 42080
rect 26160 42050 26190 42080
rect 21880 41810 21910 41850
rect 22120 41810 22150 41850
rect 22360 41810 22390 41850
rect 22600 41810 22630 41850
rect 22840 41810 22870 41850
rect 23080 41810 23110 41850
rect 23320 41810 23350 41850
rect 23560 41810 23590 41850
rect 23880 41810 23910 41850
rect 24480 41810 24510 41850
rect 24720 41810 24750 41850
rect 24960 41810 24990 41850
rect 25200 41810 25230 41850
rect 25440 41810 25470 41850
rect 25680 41810 25710 41850
rect 25920 41810 25950 41850
rect 26160 41810 26190 41850
rect 21880 41800 21990 41810
rect 21880 41760 21930 41800
rect 21970 41760 21990 41800
rect 21880 41750 21990 41760
rect 22120 41800 22230 41810
rect 22120 41760 22170 41800
rect 22210 41760 22230 41800
rect 22120 41750 22230 41760
rect 22360 41800 22470 41810
rect 22360 41760 22410 41800
rect 22450 41760 22470 41800
rect 22360 41750 22470 41760
rect 22600 41800 22710 41810
rect 22600 41760 22650 41800
rect 22690 41760 22710 41800
rect 22600 41750 22710 41760
rect 22840 41800 22950 41810
rect 22840 41760 22890 41800
rect 22930 41760 22950 41800
rect 22840 41750 22950 41760
rect 23080 41800 23190 41810
rect 23080 41760 23130 41800
rect 23170 41760 23190 41800
rect 23080 41750 23190 41760
rect 23320 41800 23430 41810
rect 23320 41760 23370 41800
rect 23410 41760 23430 41800
rect 23320 41750 23430 41760
rect 23560 41800 23670 41810
rect 23560 41760 23610 41800
rect 23650 41760 23670 41800
rect 23560 41750 23670 41760
rect 23770 41800 23910 41810
rect 23770 41720 23790 41800
rect 23870 41720 23910 41800
rect 24410 41800 24510 41810
rect 24410 41760 24430 41800
rect 24470 41760 24510 41800
rect 24410 41750 24510 41760
rect 24650 41800 24750 41810
rect 24650 41760 24670 41800
rect 24710 41760 24750 41800
rect 24650 41750 24750 41760
rect 24890 41800 24990 41810
rect 24890 41760 24910 41800
rect 24950 41760 24990 41800
rect 24890 41750 24990 41760
rect 25130 41800 25230 41810
rect 25130 41760 25150 41800
rect 25190 41760 25230 41800
rect 25130 41750 25230 41760
rect 25370 41800 25470 41810
rect 25370 41760 25390 41800
rect 25430 41760 25470 41800
rect 25370 41750 25470 41760
rect 25610 41800 25710 41810
rect 25610 41760 25630 41800
rect 25670 41760 25710 41800
rect 25610 41750 25710 41760
rect 25850 41800 25950 41810
rect 25850 41760 25870 41800
rect 25910 41760 25950 41800
rect 25850 41750 25950 41760
rect 26090 41800 26190 41810
rect 26090 41760 26110 41800
rect 26150 41760 26190 41800
rect 26090 41750 26190 41760
rect 23770 41710 23910 41720
rect 24200 41720 24330 41730
rect 21810 41690 21910 41700
rect 21810 41650 21830 41690
rect 21870 41650 21910 41690
rect 21810 41640 21910 41650
rect 22050 41690 22150 41700
rect 22050 41650 22070 41690
rect 22110 41650 22150 41690
rect 22050 41640 22150 41650
rect 22290 41690 22390 41700
rect 22290 41650 22310 41690
rect 22350 41650 22390 41690
rect 22290 41640 22390 41650
rect 22530 41690 22630 41700
rect 22530 41650 22550 41690
rect 22590 41650 22630 41690
rect 22530 41640 22630 41650
rect 22770 41690 22870 41700
rect 22770 41650 22790 41690
rect 22830 41650 22870 41690
rect 22770 41640 22870 41650
rect 23010 41690 23110 41700
rect 23010 41650 23030 41690
rect 23070 41650 23110 41690
rect 23010 41640 23110 41650
rect 23250 41690 23350 41700
rect 23250 41650 23270 41690
rect 23310 41650 23350 41690
rect 23250 41640 23350 41650
rect 23490 41690 23590 41700
rect 23490 41650 23510 41690
rect 23550 41650 23590 41690
rect 23490 41640 23590 41650
rect 21880 41604 21910 41640
rect 22120 41604 22150 41640
rect 22360 41604 22390 41640
rect 22600 41604 22630 41640
rect 22840 41604 22870 41640
rect 23080 41604 23110 41640
rect 23320 41604 23350 41640
rect 23560 41604 23590 41640
rect 24200 41650 24240 41720
rect 24310 41650 24330 41720
rect 24200 41640 24330 41650
rect 24480 41690 24570 41700
rect 24480 41650 24510 41690
rect 24550 41650 24570 41690
rect 24480 41640 24570 41650
rect 24720 41690 24810 41700
rect 24720 41650 24750 41690
rect 24790 41650 24810 41690
rect 24720 41640 24810 41650
rect 24960 41690 25050 41700
rect 24960 41650 24990 41690
rect 25030 41650 25050 41690
rect 24960 41640 25050 41650
rect 25200 41690 25290 41700
rect 25200 41650 25230 41690
rect 25270 41650 25290 41690
rect 25200 41640 25290 41650
rect 25440 41690 25530 41700
rect 25440 41650 25470 41690
rect 25510 41650 25530 41690
rect 25440 41640 25530 41650
rect 25680 41690 25770 41700
rect 25680 41650 25710 41690
rect 25750 41650 25770 41690
rect 25680 41640 25770 41650
rect 25920 41690 26010 41700
rect 25920 41650 25950 41690
rect 25990 41650 26010 41690
rect 25920 41640 26010 41650
rect 26160 41690 26250 41700
rect 26160 41650 26190 41690
rect 26230 41650 26250 41690
rect 26160 41640 26250 41650
rect 24200 41604 24230 41640
rect 24480 41604 24510 41640
rect 24720 41604 24750 41640
rect 24960 41604 24990 41640
rect 25200 41604 25230 41640
rect 25440 41604 25470 41640
rect 25680 41604 25710 41640
rect 25920 41604 25950 41640
rect 26160 41604 26190 41640
rect 21880 41490 21910 41520
rect 22120 41490 22150 41520
rect 22360 41490 22390 41520
rect 22600 41490 22630 41520
rect 22840 41490 22870 41520
rect 23080 41490 23110 41520
rect 23320 41490 23350 41520
rect 23560 41490 23590 41520
rect 24200 41490 24230 41520
rect 24480 41490 24510 41520
rect 24720 41490 24750 41520
rect 24960 41490 24990 41520
rect 25200 41490 25230 41520
rect 25440 41490 25470 41520
rect 25680 41490 25710 41520
rect 25920 41490 25950 41520
rect 26160 41490 26190 41520
rect 23810 41210 23840 41240
rect 24140 41210 24170 41240
rect 24400 41210 24430 41240
rect 23810 40890 23840 41010
rect 24140 40970 24170 41010
rect 24400 40970 24430 41010
rect 24060 40960 24170 40970
rect 24060 40920 24080 40960
rect 24120 40920 24170 40960
rect 24060 40910 24170 40920
rect 24320 40960 24430 40970
rect 24320 40920 24340 40960
rect 24380 40920 24430 40960
rect 24320 40910 24430 40920
rect 23810 40880 24020 40890
rect 23810 40840 23960 40880
rect 24000 40840 24020 40880
rect 23810 40830 24020 40840
rect 23810 40794 23840 40830
rect 24140 40794 24170 40910
rect 24400 40794 24430 40910
rect 23810 40680 23840 40710
rect 24140 40680 24170 40710
rect 24400 40680 24430 40710
rect 21880 39460 21910 39490
rect 22120 39460 22150 39490
rect 22360 39460 22390 39490
rect 22600 39460 22630 39490
rect 22840 39460 22870 39490
rect 23080 39460 23110 39490
rect 23320 39460 23350 39490
rect 23560 39460 23590 39490
rect 23880 39460 23910 39490
rect 24480 39460 24510 39490
rect 24720 39460 24750 39490
rect 24960 39460 24990 39490
rect 25200 39460 25230 39490
rect 25440 39460 25470 39490
rect 25680 39460 25710 39490
rect 25920 39460 25950 39490
rect 26160 39460 26190 39490
rect 13070 39210 13100 39240
rect 13400 39210 13430 39240
rect 21880 39220 21910 39260
rect 22120 39220 22150 39260
rect 22360 39220 22390 39260
rect 22600 39220 22630 39260
rect 22840 39220 22870 39260
rect 23080 39220 23110 39260
rect 23320 39220 23350 39260
rect 23560 39220 23590 39260
rect 23880 39220 23910 39260
rect 24480 39220 24510 39260
rect 24720 39220 24750 39260
rect 24960 39220 24990 39260
rect 25200 39220 25230 39260
rect 25440 39220 25470 39260
rect 25680 39220 25710 39260
rect 25920 39220 25950 39260
rect 26160 39220 26190 39260
rect 21880 39210 21990 39220
rect 21880 39170 21930 39210
rect 21970 39170 21990 39210
rect 21880 39160 21990 39170
rect 22120 39210 22230 39220
rect 22120 39170 22170 39210
rect 22210 39170 22230 39210
rect 22120 39160 22230 39170
rect 22360 39210 22470 39220
rect 22360 39170 22410 39210
rect 22450 39170 22470 39210
rect 22360 39160 22470 39170
rect 22600 39210 22710 39220
rect 22600 39170 22650 39210
rect 22690 39170 22710 39210
rect 22600 39160 22710 39170
rect 22840 39210 22950 39220
rect 22840 39170 22890 39210
rect 22930 39170 22950 39210
rect 22840 39160 22950 39170
rect 23080 39210 23190 39220
rect 23080 39170 23130 39210
rect 23170 39170 23190 39210
rect 23080 39160 23190 39170
rect 23320 39210 23430 39220
rect 23320 39170 23370 39210
rect 23410 39170 23430 39210
rect 23320 39160 23430 39170
rect 23560 39210 23670 39220
rect 23560 39170 23610 39210
rect 23650 39170 23670 39210
rect 23560 39160 23670 39170
rect 23770 39210 23910 39220
rect 23770 39130 23790 39210
rect 23870 39130 23910 39210
rect 24410 39210 24510 39220
rect 24410 39170 24430 39210
rect 24470 39170 24510 39210
rect 24410 39160 24510 39170
rect 24650 39210 24750 39220
rect 24650 39170 24670 39210
rect 24710 39170 24750 39210
rect 24650 39160 24750 39170
rect 24890 39210 24990 39220
rect 24890 39170 24910 39210
rect 24950 39170 24990 39210
rect 24890 39160 24990 39170
rect 25130 39210 25230 39220
rect 25130 39170 25150 39210
rect 25190 39170 25230 39210
rect 25130 39160 25230 39170
rect 25370 39210 25470 39220
rect 25370 39170 25390 39210
rect 25430 39170 25470 39210
rect 25370 39160 25470 39170
rect 25610 39210 25710 39220
rect 25610 39170 25630 39210
rect 25670 39170 25710 39210
rect 25610 39160 25710 39170
rect 25850 39210 25950 39220
rect 25850 39170 25870 39210
rect 25910 39170 25950 39210
rect 25850 39160 25950 39170
rect 26090 39210 26190 39220
rect 26090 39170 26110 39210
rect 26150 39170 26190 39210
rect 26090 39160 26190 39170
rect 23770 39120 23910 39130
rect 24200 39130 24330 39140
rect 21810 39100 21910 39110
rect 21810 39060 21830 39100
rect 21870 39060 21910 39100
rect 21810 39050 21910 39060
rect 22050 39100 22150 39110
rect 22050 39060 22070 39100
rect 22110 39060 22150 39100
rect 22050 39050 22150 39060
rect 22290 39100 22390 39110
rect 22290 39060 22310 39100
rect 22350 39060 22390 39100
rect 22290 39050 22390 39060
rect 22530 39100 22630 39110
rect 22530 39060 22550 39100
rect 22590 39060 22630 39100
rect 22530 39050 22630 39060
rect 22770 39100 22870 39110
rect 22770 39060 22790 39100
rect 22830 39060 22870 39100
rect 22770 39050 22870 39060
rect 23010 39100 23110 39110
rect 23010 39060 23030 39100
rect 23070 39060 23110 39100
rect 23010 39050 23110 39060
rect 23250 39100 23350 39110
rect 23250 39060 23270 39100
rect 23310 39060 23350 39100
rect 23250 39050 23350 39060
rect 23490 39100 23590 39110
rect 23490 39060 23510 39100
rect 23550 39060 23590 39100
rect 23490 39050 23590 39060
rect 21880 39014 21910 39050
rect 22120 39014 22150 39050
rect 22360 39014 22390 39050
rect 22600 39014 22630 39050
rect 22840 39014 22870 39050
rect 23080 39014 23110 39050
rect 23320 39014 23350 39050
rect 23560 39014 23590 39050
rect 24200 39060 24240 39130
rect 24310 39060 24330 39130
rect 24200 39050 24330 39060
rect 24480 39100 24570 39110
rect 24480 39060 24510 39100
rect 24550 39060 24570 39100
rect 24480 39050 24570 39060
rect 24720 39100 24810 39110
rect 24720 39060 24750 39100
rect 24790 39060 24810 39100
rect 24720 39050 24810 39060
rect 24960 39100 25050 39110
rect 24960 39060 24990 39100
rect 25030 39060 25050 39100
rect 24960 39050 25050 39060
rect 25200 39100 25290 39110
rect 25200 39060 25230 39100
rect 25270 39060 25290 39100
rect 25200 39050 25290 39060
rect 25440 39100 25530 39110
rect 25440 39060 25470 39100
rect 25510 39060 25530 39100
rect 25440 39050 25530 39060
rect 25680 39100 25770 39110
rect 25680 39060 25710 39100
rect 25750 39060 25770 39100
rect 25680 39050 25770 39060
rect 25920 39100 26010 39110
rect 25920 39060 25950 39100
rect 25990 39060 26010 39100
rect 25920 39050 26010 39060
rect 26160 39100 26250 39110
rect 26160 39060 26190 39100
rect 26230 39060 26250 39100
rect 26160 39050 26250 39060
rect 24200 39014 24230 39050
rect 24480 39014 24510 39050
rect 24720 39014 24750 39050
rect 24960 39014 24990 39050
rect 25200 39014 25230 39050
rect 25440 39014 25470 39050
rect 25680 39014 25710 39050
rect 25920 39014 25950 39050
rect 26160 39014 26190 39050
rect 13070 38890 13100 39010
rect 13400 38970 13430 39010
rect 13320 38960 13430 38970
rect 13320 38920 13340 38960
rect 13380 38920 13430 38960
rect 13320 38910 13430 38920
rect 13070 38880 13280 38890
rect 13070 38840 13220 38880
rect 13260 38840 13280 38880
rect 13070 38830 13280 38840
rect 13070 38794 13100 38830
rect 13400 38794 13430 38910
rect 21880 38900 21910 38930
rect 22120 38900 22150 38930
rect 22360 38900 22390 38930
rect 22600 38900 22630 38930
rect 22840 38900 22870 38930
rect 23080 38900 23110 38930
rect 23320 38900 23350 38930
rect 23560 38900 23590 38930
rect 24200 38900 24230 38930
rect 24480 38900 24510 38930
rect 24720 38900 24750 38930
rect 24960 38900 24990 38930
rect 25200 38900 25230 38930
rect 25440 38900 25470 38930
rect 25680 38900 25710 38930
rect 25920 38900 25950 38930
rect 26160 38900 26190 38930
rect 13070 38680 13100 38710
rect 13400 38680 13430 38710
<< polycont >>
rect 21930 41760 21970 41800
rect 22170 41760 22210 41800
rect 22410 41760 22450 41800
rect 22650 41760 22690 41800
rect 22890 41760 22930 41800
rect 23130 41760 23170 41800
rect 23370 41760 23410 41800
rect 23610 41760 23650 41800
rect 23790 41720 23870 41800
rect 24430 41760 24470 41800
rect 24670 41760 24710 41800
rect 24910 41760 24950 41800
rect 25150 41760 25190 41800
rect 25390 41760 25430 41800
rect 25630 41760 25670 41800
rect 25870 41760 25910 41800
rect 26110 41760 26150 41800
rect 21830 41650 21870 41690
rect 22070 41650 22110 41690
rect 22310 41650 22350 41690
rect 22550 41650 22590 41690
rect 22790 41650 22830 41690
rect 23030 41650 23070 41690
rect 23270 41650 23310 41690
rect 23510 41650 23550 41690
rect 24240 41650 24310 41720
rect 24510 41650 24550 41690
rect 24750 41650 24790 41690
rect 24990 41650 25030 41690
rect 25230 41650 25270 41690
rect 25470 41650 25510 41690
rect 25710 41650 25750 41690
rect 25950 41650 25990 41690
rect 26190 41650 26230 41690
rect 24080 40920 24120 40960
rect 24340 40920 24380 40960
rect 23960 40840 24000 40880
rect 21930 39170 21970 39210
rect 22170 39170 22210 39210
rect 22410 39170 22450 39210
rect 22650 39170 22690 39210
rect 22890 39170 22930 39210
rect 23130 39170 23170 39210
rect 23370 39170 23410 39210
rect 23610 39170 23650 39210
rect 23790 39130 23870 39210
rect 24430 39170 24470 39210
rect 24670 39170 24710 39210
rect 24910 39170 24950 39210
rect 25150 39170 25190 39210
rect 25390 39170 25430 39210
rect 25630 39170 25670 39210
rect 25870 39170 25910 39210
rect 26110 39170 26150 39210
rect 21830 39060 21870 39100
rect 22070 39060 22110 39100
rect 22310 39060 22350 39100
rect 22550 39060 22590 39100
rect 22790 39060 22830 39100
rect 23030 39060 23070 39100
rect 23270 39060 23310 39100
rect 23510 39060 23550 39100
rect 24240 39060 24310 39130
rect 24510 39060 24550 39100
rect 24750 39060 24790 39100
rect 24990 39060 25030 39100
rect 25230 39060 25270 39100
rect 25470 39060 25510 39100
rect 25710 39060 25750 39100
rect 25950 39060 25990 39100
rect 26190 39060 26230 39100
rect 13340 38920 13380 38960
rect 13220 38840 13260 38880
<< locali >>
rect 21140 42150 26790 42170
rect 21140 42110 21160 42150
rect 21200 42110 21730 42150
rect 21770 42110 21890 42150
rect 21930 42110 22050 42150
rect 22090 42110 22210 42150
rect 22250 42110 22370 42150
rect 22410 42110 22530 42150
rect 22570 42110 22690 42150
rect 22730 42110 22850 42150
rect 22890 42110 23010 42150
rect 23050 42110 23170 42150
rect 23210 42110 23330 42150
rect 23370 42110 23490 42150
rect 23530 42110 23650 42150
rect 23690 42110 23810 42150
rect 23850 42110 23970 42150
rect 24010 42110 24330 42150
rect 24370 42110 24490 42150
rect 24530 42110 24650 42150
rect 24690 42110 24810 42150
rect 24850 42110 24970 42150
rect 25010 42110 25130 42150
rect 25170 42110 25290 42150
rect 25330 42110 25450 42150
rect 25490 42110 25610 42150
rect 25650 42110 25770 42150
rect 25810 42110 25930 42150
rect 25970 42110 26090 42150
rect 26130 42110 26250 42150
rect 26290 42110 26730 42150
rect 26770 42110 26790 42150
rect 21140 42090 26790 42110
rect 21800 42020 21860 42090
rect 21800 41880 21820 42020
rect 21800 41850 21860 41880
rect 21930 42020 21970 42050
rect 21930 41810 21970 41880
rect 22040 42020 22100 42090
rect 22040 41880 22060 42020
rect 22040 41850 22100 41880
rect 22170 42020 22210 42050
rect 22170 41810 22210 41880
rect 22280 42020 22340 42090
rect 22280 41880 22300 42020
rect 22280 41850 22340 41880
rect 22410 42020 22450 42050
rect 22410 41810 22450 41880
rect 22520 42020 22580 42090
rect 22520 41880 22540 42020
rect 22520 41850 22580 41880
rect 22650 42020 22690 42050
rect 22650 41810 22690 41880
rect 22760 42020 22820 42090
rect 22760 41880 22780 42020
rect 22760 41850 22820 41880
rect 22890 42020 22930 42050
rect 22890 41810 22930 41880
rect 23000 42020 23060 42090
rect 23000 41880 23020 42020
rect 23000 41850 23060 41880
rect 23130 42020 23170 42050
rect 23130 41810 23170 41880
rect 23240 42020 23300 42090
rect 23240 41880 23260 42020
rect 23240 41850 23300 41880
rect 23370 42020 23410 42050
rect 23370 41810 23410 41880
rect 23480 42020 23540 42090
rect 23480 41880 23500 42020
rect 23480 41850 23540 41880
rect 23610 42020 23650 42050
rect 23610 41810 23650 41880
rect 23780 42020 23860 42090
rect 23780 41850 23860 41880
rect 23930 42020 24010 42050
rect 21780 41800 23890 41810
rect 21780 41760 21930 41800
rect 21970 41760 22170 41800
rect 22210 41760 22410 41800
rect 22450 41760 22650 41800
rect 22690 41760 22890 41800
rect 22930 41760 23130 41800
rect 23170 41760 23370 41800
rect 23410 41760 23610 41800
rect 23650 41760 23790 41800
rect 21780 41730 23790 41760
rect 21150 41660 21550 41680
rect 21150 41620 21170 41660
rect 21210 41620 21550 41660
rect 21810 41650 21830 41690
rect 21870 41650 21890 41690
rect 21150 41600 21550 41620
rect 21470 41480 21550 41600
rect 21800 41580 21860 41600
rect 21800 41540 21820 41580
rect 21800 41480 21860 41540
rect 21930 41580 21970 41730
rect 22050 41650 22070 41690
rect 22110 41650 22130 41690
rect 21930 41520 21970 41540
rect 22040 41580 22100 41600
rect 22040 41540 22060 41580
rect 22040 41480 22100 41540
rect 22170 41580 22210 41730
rect 22290 41650 22310 41690
rect 22350 41650 22370 41690
rect 22170 41520 22210 41540
rect 22280 41580 22340 41600
rect 22280 41540 22300 41580
rect 22280 41480 22340 41540
rect 22410 41580 22450 41730
rect 22530 41650 22550 41690
rect 22590 41650 22610 41690
rect 22410 41520 22450 41540
rect 22520 41580 22580 41600
rect 22520 41540 22540 41580
rect 22520 41480 22580 41540
rect 22650 41580 22690 41730
rect 22770 41650 22790 41690
rect 22830 41650 22850 41690
rect 22650 41520 22690 41540
rect 22760 41580 22820 41600
rect 22760 41540 22780 41580
rect 22760 41480 22820 41540
rect 22890 41580 22930 41730
rect 23010 41650 23030 41690
rect 23070 41650 23090 41690
rect 22890 41520 22930 41540
rect 23000 41580 23060 41600
rect 23000 41540 23020 41580
rect 23000 41480 23060 41540
rect 23130 41580 23170 41730
rect 23250 41650 23270 41690
rect 23310 41650 23330 41690
rect 23130 41520 23170 41540
rect 23240 41580 23300 41600
rect 23240 41540 23260 41580
rect 23240 41480 23300 41540
rect 23370 41580 23410 41730
rect 23610 41720 23790 41730
rect 23870 41720 23890 41800
rect 23610 41710 23890 41720
rect 23490 41650 23510 41690
rect 23550 41650 23570 41690
rect 23370 41520 23410 41540
rect 23480 41580 23540 41600
rect 23480 41540 23500 41580
rect 23480 41480 23540 41540
rect 23610 41580 23650 41710
rect 23610 41520 23650 41540
rect 23930 41600 24010 41880
rect 24400 42020 24460 42090
rect 24400 41880 24420 42020
rect 24400 41850 24460 41880
rect 24530 42020 24570 42050
rect 24410 41800 24490 41810
rect 24410 41760 24430 41800
rect 24470 41760 24490 41800
rect 24410 41750 24490 41760
rect 24220 41720 24330 41730
rect 24220 41650 24240 41720
rect 24310 41710 24330 41720
rect 24530 41710 24570 41880
rect 24640 42020 24700 42090
rect 24640 41880 24660 42020
rect 24640 41850 24700 41880
rect 24770 42020 24810 42050
rect 24650 41800 24730 41810
rect 24650 41760 24670 41800
rect 24710 41760 24730 41800
rect 24650 41750 24730 41760
rect 24770 41710 24810 41880
rect 24880 42020 24940 42090
rect 24880 41880 24900 42020
rect 24880 41850 24940 41880
rect 25010 42020 25050 42050
rect 24890 41800 24970 41810
rect 24890 41760 24910 41800
rect 24950 41760 24970 41800
rect 24890 41750 24970 41760
rect 25010 41710 25050 41880
rect 25120 42020 25180 42090
rect 25120 41880 25140 42020
rect 25120 41850 25180 41880
rect 25250 42020 25290 42050
rect 25130 41800 25210 41810
rect 25130 41760 25150 41800
rect 25190 41760 25210 41800
rect 25130 41750 25210 41760
rect 25250 41710 25290 41880
rect 25360 42020 25420 42090
rect 25360 41880 25380 42020
rect 25360 41850 25420 41880
rect 25490 42020 25530 42050
rect 25370 41800 25450 41810
rect 25370 41760 25390 41800
rect 25430 41760 25450 41800
rect 25370 41750 25450 41760
rect 25490 41710 25530 41880
rect 25600 42020 25660 42090
rect 25600 41880 25620 42020
rect 25600 41850 25660 41880
rect 25730 42020 25770 42050
rect 25610 41800 25690 41810
rect 25610 41760 25630 41800
rect 25670 41760 25690 41800
rect 25610 41750 25690 41760
rect 25730 41710 25770 41880
rect 25840 42020 25900 42090
rect 25840 41880 25860 42020
rect 25840 41850 25900 41880
rect 25970 42020 26010 42050
rect 25850 41800 25930 41810
rect 25850 41760 25870 41800
rect 25910 41760 25930 41800
rect 25850 41750 25930 41760
rect 25970 41710 26010 41880
rect 26080 42020 26140 42090
rect 26080 41880 26100 42020
rect 26080 41850 26140 41880
rect 26210 42020 26250 42050
rect 26090 41800 26170 41810
rect 26090 41760 26110 41800
rect 26150 41760 26170 41800
rect 26090 41750 26170 41760
rect 26210 41710 26250 41880
rect 24310 41690 26250 41710
rect 24310 41650 24510 41690
rect 24550 41650 24750 41690
rect 24790 41650 24990 41690
rect 25030 41650 25230 41690
rect 25270 41650 25470 41690
rect 25510 41650 25710 41690
rect 25750 41650 25950 41690
rect 25990 41650 26190 41690
rect 26230 41650 26250 41690
rect 24220 41640 26250 41650
rect 23930 41580 24180 41600
rect 23930 41540 23950 41580
rect 23990 41540 24100 41580
rect 23930 41520 24180 41540
rect 24250 41580 24330 41600
rect 24250 41480 24330 41540
rect 24420 41580 24460 41600
rect 24420 41480 24460 41540
rect 24530 41580 24570 41640
rect 24530 41520 24570 41540
rect 24640 41580 24700 41600
rect 24640 41540 24660 41580
rect 24640 41480 24700 41540
rect 24770 41580 24810 41640
rect 24770 41520 24810 41540
rect 24900 41580 24940 41600
rect 24900 41480 24940 41540
rect 25010 41580 25050 41640
rect 25010 41520 25050 41540
rect 25120 41580 25180 41600
rect 25120 41540 25140 41580
rect 25120 41480 25180 41540
rect 25250 41580 25290 41640
rect 25250 41520 25290 41540
rect 25380 41580 25420 41600
rect 25380 41480 25420 41540
rect 25490 41580 25530 41640
rect 25490 41520 25530 41540
rect 25600 41580 25660 41600
rect 25600 41540 25620 41580
rect 25600 41480 25660 41540
rect 25730 41580 25770 41640
rect 25730 41520 25770 41540
rect 25860 41580 25900 41600
rect 25860 41480 25900 41540
rect 25970 41580 26010 41640
rect 25970 41520 26010 41540
rect 26080 41580 26140 41600
rect 26080 41540 26100 41580
rect 26080 41480 26140 41540
rect 26210 41580 26250 41640
rect 26210 41520 26250 41540
rect 21470 41460 26540 41480
rect 21470 41420 21730 41460
rect 21770 41420 21890 41460
rect 21930 41420 22050 41460
rect 22090 41420 22210 41460
rect 22250 41420 22370 41460
rect 22410 41420 22530 41460
rect 22570 41420 22690 41460
rect 22730 41420 22850 41460
rect 22890 41420 23010 41460
rect 23050 41420 23170 41460
rect 23210 41420 23330 41460
rect 23370 41420 23490 41460
rect 23530 41420 23650 41460
rect 23690 41420 24170 41460
rect 24210 41420 24330 41460
rect 24370 41420 24490 41460
rect 24530 41420 24650 41460
rect 24690 41420 24810 41460
rect 24850 41420 24970 41460
rect 25010 41420 25130 41460
rect 25170 41420 25290 41460
rect 25330 41420 25450 41460
rect 25490 41420 25610 41460
rect 25650 41420 25770 41460
rect 25810 41420 25930 41460
rect 25970 41420 26090 41460
rect 26130 41420 26250 41460
rect 26290 41420 26540 41460
rect 21470 41400 26540 41420
rect 21140 41310 26340 41330
rect 21140 41270 21160 41310
rect 21200 41270 23750 41310
rect 23790 41270 23910 41310
rect 23950 41270 24070 41310
rect 24110 41270 24230 41310
rect 24270 41270 24390 41310
rect 24430 41270 24550 41310
rect 24590 41270 26280 41310
rect 26320 41270 26340 41310
rect 21140 41250 26340 41270
rect 23670 41180 23710 41210
rect 23670 40670 23710 41040
rect 23750 40770 23790 41250
rect 23750 40710 23790 40730
rect 23860 41180 23900 41210
rect 23860 40960 23900 41040
rect 24060 41180 24120 41250
rect 24060 41040 24080 41180
rect 24060 41010 24120 41040
rect 24190 41180 24250 41210
rect 24230 41040 24250 41180
rect 24190 40960 24250 41040
rect 24320 41180 24380 41250
rect 24320 41040 24340 41180
rect 24320 41010 24380 41040
rect 24450 41180 24510 41210
rect 24490 41040 24510 41180
rect 23860 40920 23950 40960
rect 23990 40920 24080 40960
rect 24120 40920 24140 40960
rect 24190 40920 24340 40960
rect 24380 40920 24400 40960
rect 24450 40920 24510 41040
rect 23860 40770 23900 40920
rect 24190 40880 24250 40920
rect 23940 40840 23960 40880
rect 24000 40840 24250 40880
rect 23860 40710 23900 40730
rect 24060 40770 24120 40790
rect 24060 40730 24080 40770
rect 24060 40670 24120 40730
rect 24190 40770 24250 40840
rect 24450 40870 26270 40920
rect 24230 40730 24250 40770
rect 24190 40710 24250 40730
rect 24320 40770 24380 40790
rect 24320 40730 24340 40770
rect 24320 40670 24380 40730
rect 24450 40770 24510 40870
rect 24490 40730 24510 40770
rect 24450 40710 24510 40730
rect 26460 40670 26540 41400
rect 21140 40660 26540 40670
rect 21140 40650 26480 40660
rect 21140 40610 21160 40650
rect 21200 40610 23750 40650
rect 23790 40610 23910 40650
rect 23950 40610 24070 40650
rect 24110 40610 24230 40650
rect 24270 40610 24390 40650
rect 24430 40610 24550 40650
rect 24590 40620 26480 40650
rect 26520 40620 26540 40660
rect 24590 40610 26540 40620
rect 21140 40590 26540 40610
rect 21140 39560 26790 39580
rect 21140 39520 21160 39560
rect 21200 39520 21730 39560
rect 21770 39520 21890 39560
rect 21930 39520 22050 39560
rect 22090 39520 22210 39560
rect 22250 39520 22370 39560
rect 22410 39520 22530 39560
rect 22570 39520 22690 39560
rect 22730 39520 22850 39560
rect 22890 39520 23010 39560
rect 23050 39520 23170 39560
rect 23210 39520 23330 39560
rect 23370 39520 23490 39560
rect 23530 39520 23650 39560
rect 23690 39520 23810 39560
rect 23850 39520 23970 39560
rect 24010 39520 24330 39560
rect 24370 39520 24490 39560
rect 24530 39520 24650 39560
rect 24690 39520 24810 39560
rect 24850 39520 24970 39560
rect 25010 39520 25130 39560
rect 25170 39520 25290 39560
rect 25330 39520 25450 39560
rect 25490 39520 25610 39560
rect 25650 39520 25770 39560
rect 25810 39520 25930 39560
rect 25970 39520 26090 39560
rect 26130 39520 26250 39560
rect 26290 39520 26730 39560
rect 26770 39520 26790 39560
rect 21140 39500 26790 39520
rect 21800 39430 21860 39500
rect 12708 39310 13550 39330
rect 12708 39270 13010 39310
rect 13050 39270 13170 39310
rect 13210 39270 13330 39310
rect 13370 39270 13490 39310
rect 13530 39270 13550 39310
rect 12708 39250 13550 39270
rect 21800 39290 21820 39430
rect 21800 39260 21860 39290
rect 21930 39430 21970 39460
rect 12930 39180 12970 39210
rect 12930 38670 12970 39040
rect 13010 38770 13050 39250
rect 13010 38710 13050 38730
rect 13120 39180 13160 39210
rect 13120 38960 13160 39040
rect 13320 39180 13380 39250
rect 21930 39220 21970 39290
rect 22040 39430 22100 39500
rect 22040 39290 22060 39430
rect 22040 39260 22100 39290
rect 22170 39430 22210 39460
rect 22170 39220 22210 39290
rect 22280 39430 22340 39500
rect 22280 39290 22300 39430
rect 22280 39260 22340 39290
rect 22410 39430 22450 39460
rect 22410 39220 22450 39290
rect 22520 39430 22580 39500
rect 22520 39290 22540 39430
rect 22520 39260 22580 39290
rect 22650 39430 22690 39460
rect 22650 39220 22690 39290
rect 22760 39430 22820 39500
rect 22760 39290 22780 39430
rect 22760 39260 22820 39290
rect 22890 39430 22930 39460
rect 22890 39220 22930 39290
rect 23000 39430 23060 39500
rect 23000 39290 23020 39430
rect 23000 39260 23060 39290
rect 23130 39430 23170 39460
rect 23130 39220 23170 39290
rect 23240 39430 23300 39500
rect 23240 39290 23260 39430
rect 23240 39260 23300 39290
rect 23370 39430 23410 39460
rect 23370 39220 23410 39290
rect 23480 39430 23540 39500
rect 23480 39290 23500 39430
rect 23480 39260 23540 39290
rect 23610 39430 23650 39460
rect 23610 39220 23650 39290
rect 23780 39430 23860 39500
rect 23780 39260 23860 39290
rect 23930 39430 24010 39460
rect 21780 39210 23890 39220
rect 13320 39040 13340 39180
rect 13320 39010 13380 39040
rect 13450 39180 13510 39210
rect 13490 39040 13510 39180
rect 21780 39170 21930 39210
rect 21970 39170 22170 39210
rect 22210 39170 22410 39210
rect 22450 39170 22650 39210
rect 22690 39170 22890 39210
rect 22930 39170 23130 39210
rect 23170 39170 23370 39210
rect 23410 39170 23610 39210
rect 23650 39170 23790 39210
rect 21780 39140 23790 39170
rect 13120 38920 13210 38960
rect 13250 38920 13340 38960
rect 13380 38920 13400 38960
rect 13450 38920 13510 39040
rect 21810 39060 21830 39100
rect 21870 39060 21890 39100
rect 14210 38920 14260 39040
rect 13120 38770 13160 38920
rect 13450 38880 13618 38920
rect 14140 38880 14260 38920
rect 21800 38990 21860 39010
rect 21800 38950 21820 38990
rect 21800 38890 21860 38950
rect 21930 38990 21970 39140
rect 22050 39060 22070 39100
rect 22110 39060 22130 39100
rect 21930 38930 21970 38950
rect 22040 38990 22100 39010
rect 22040 38950 22060 38990
rect 22040 38890 22100 38950
rect 22170 38990 22210 39140
rect 22290 39060 22310 39100
rect 22350 39060 22370 39100
rect 22170 38930 22210 38950
rect 22280 38990 22340 39010
rect 22280 38950 22300 38990
rect 22280 38890 22340 38950
rect 22410 38990 22450 39140
rect 22530 39060 22550 39100
rect 22590 39060 22610 39100
rect 22410 38930 22450 38950
rect 22520 38990 22580 39010
rect 22520 38950 22540 38990
rect 22520 38890 22580 38950
rect 22650 38990 22690 39140
rect 22770 39060 22790 39100
rect 22830 39060 22850 39100
rect 22650 38930 22690 38950
rect 22760 38990 22820 39010
rect 22760 38950 22780 38990
rect 22760 38890 22820 38950
rect 22890 38990 22930 39140
rect 23010 39060 23030 39100
rect 23070 39060 23090 39100
rect 22890 38930 22930 38950
rect 23000 38990 23060 39010
rect 23000 38950 23020 38990
rect 23000 38890 23060 38950
rect 23130 38990 23170 39140
rect 23250 39060 23270 39100
rect 23310 39060 23330 39100
rect 23130 38930 23170 38950
rect 23240 38990 23300 39010
rect 23240 38950 23260 38990
rect 23240 38890 23300 38950
rect 23370 38990 23410 39140
rect 23610 39130 23790 39140
rect 23870 39130 23890 39210
rect 23610 39120 23890 39130
rect 23490 39060 23510 39100
rect 23550 39060 23570 39100
rect 23370 38930 23410 38950
rect 23480 38990 23540 39010
rect 23480 38950 23500 38990
rect 23480 38890 23540 38950
rect 23610 38990 23650 39120
rect 23610 38930 23650 38950
rect 23930 39010 24010 39290
rect 24400 39430 24460 39500
rect 24400 39290 24420 39430
rect 24400 39260 24460 39290
rect 24530 39430 24570 39460
rect 24410 39210 24490 39220
rect 24410 39170 24430 39210
rect 24470 39170 24490 39210
rect 24410 39160 24490 39170
rect 24220 39130 24330 39140
rect 24220 39060 24240 39130
rect 24310 39120 24330 39130
rect 24530 39120 24570 39290
rect 24640 39430 24700 39500
rect 24640 39290 24660 39430
rect 24640 39260 24700 39290
rect 24770 39430 24810 39460
rect 24650 39210 24730 39220
rect 24650 39170 24670 39210
rect 24710 39170 24730 39210
rect 24650 39160 24730 39170
rect 24770 39120 24810 39290
rect 24880 39430 24940 39500
rect 24880 39290 24900 39430
rect 24880 39260 24940 39290
rect 25010 39430 25050 39460
rect 24890 39210 24970 39220
rect 24890 39170 24910 39210
rect 24950 39170 24970 39210
rect 24890 39160 24970 39170
rect 25010 39120 25050 39290
rect 25120 39430 25180 39500
rect 25120 39290 25140 39430
rect 25120 39260 25180 39290
rect 25250 39430 25290 39460
rect 25130 39210 25210 39220
rect 25130 39170 25150 39210
rect 25190 39170 25210 39210
rect 25130 39160 25210 39170
rect 25250 39120 25290 39290
rect 25360 39430 25420 39500
rect 25360 39290 25380 39430
rect 25360 39260 25420 39290
rect 25490 39430 25530 39460
rect 25370 39210 25450 39220
rect 25370 39170 25390 39210
rect 25430 39170 25450 39210
rect 25370 39160 25450 39170
rect 25490 39120 25530 39290
rect 25600 39430 25660 39500
rect 25600 39290 25620 39430
rect 25600 39260 25660 39290
rect 25730 39430 25770 39460
rect 25610 39210 25690 39220
rect 25610 39170 25630 39210
rect 25670 39170 25690 39210
rect 25610 39160 25690 39170
rect 25730 39120 25770 39290
rect 25840 39430 25900 39500
rect 25840 39290 25860 39430
rect 25840 39260 25900 39290
rect 25970 39430 26010 39460
rect 25850 39210 25930 39220
rect 25850 39170 25870 39210
rect 25910 39170 25930 39210
rect 25850 39160 25930 39170
rect 25970 39120 26010 39290
rect 26080 39430 26140 39500
rect 26080 39290 26100 39430
rect 26080 39260 26140 39290
rect 26210 39430 26250 39460
rect 26090 39210 26170 39220
rect 26090 39170 26110 39210
rect 26150 39170 26170 39210
rect 26090 39160 26170 39170
rect 26210 39120 26250 39290
rect 24310 39100 26250 39120
rect 24310 39060 24510 39100
rect 24550 39060 24750 39100
rect 24790 39060 24990 39100
rect 25030 39060 25230 39100
rect 25270 39060 25470 39100
rect 25510 39060 25710 39100
rect 25750 39060 25950 39100
rect 25990 39060 26190 39100
rect 26230 39060 26250 39100
rect 24220 39050 26250 39060
rect 23930 38990 24180 39010
rect 23930 38950 23950 38990
rect 23990 38950 24100 38990
rect 23930 38930 24180 38950
rect 24250 38990 24330 39010
rect 24250 38890 24330 38950
rect 24420 38990 24460 39010
rect 24420 38890 24460 38950
rect 24530 38990 24570 39050
rect 24530 38930 24570 38950
rect 24640 38990 24700 39010
rect 24640 38950 24660 38990
rect 24640 38890 24700 38950
rect 24770 38990 24810 39050
rect 24770 38930 24810 38950
rect 24900 38990 24940 39010
rect 24900 38890 24940 38950
rect 25010 38990 25050 39050
rect 25010 38930 25050 38950
rect 25120 38990 25180 39010
rect 25120 38950 25140 38990
rect 25120 38890 25180 38950
rect 25250 38990 25290 39050
rect 25250 38930 25290 38950
rect 25380 38990 25420 39010
rect 25380 38890 25420 38950
rect 25490 38990 25530 39050
rect 25490 38930 25530 38950
rect 25600 38990 25660 39010
rect 25600 38950 25620 38990
rect 25600 38890 25660 38950
rect 25730 38990 25770 39050
rect 25730 38930 25770 38950
rect 25860 38990 25900 39010
rect 25860 38890 25900 38950
rect 25970 38990 26010 39050
rect 25970 38930 26010 38950
rect 26080 38990 26140 39010
rect 26080 38950 26100 38990
rect 26080 38890 26140 38950
rect 26210 38990 26250 39050
rect 26210 38930 26250 38950
rect 21140 38880 26540 38890
rect 13200 38840 13220 38880
rect 13260 38840 13510 38880
rect 13120 38710 13160 38730
rect 13320 38770 13380 38790
rect 13320 38730 13340 38770
rect 13320 38670 13380 38730
rect 13450 38770 13510 38840
rect 21140 38870 26480 38880
rect 21140 38830 21160 38870
rect 21200 38830 21730 38870
rect 21770 38830 21890 38870
rect 21930 38830 22050 38870
rect 22090 38830 22210 38870
rect 22250 38830 22370 38870
rect 22410 38830 22530 38870
rect 22570 38830 22690 38870
rect 22730 38830 22850 38870
rect 22890 38830 23010 38870
rect 23050 38830 23170 38870
rect 23210 38830 23330 38870
rect 23370 38830 23490 38870
rect 23530 38830 23650 38870
rect 23690 38830 24170 38870
rect 24210 38830 24330 38870
rect 24370 38830 24490 38870
rect 24530 38830 24650 38870
rect 24690 38830 24810 38870
rect 24850 38830 24970 38870
rect 25010 38830 25130 38870
rect 25170 38830 25290 38870
rect 25330 38830 25450 38870
rect 25490 38830 25610 38870
rect 25650 38830 25770 38870
rect 25810 38830 25930 38870
rect 25970 38830 26090 38870
rect 26130 38830 26250 38870
rect 26290 38840 26480 38870
rect 26520 38840 26540 38880
rect 26290 38830 26540 38840
rect 21140 38810 26540 38830
rect 13490 38730 13510 38770
rect 13450 38710 13510 38730
rect 12708 38650 13550 38670
rect 12708 38610 13010 38650
rect 13050 38610 13170 38650
rect 13210 38610 13330 38650
rect 13370 38610 13490 38650
rect 13530 38610 13550 38650
rect 12708 38590 13550 38610
<< viali >>
rect 21160 42110 21200 42150
rect 26730 42110 26770 42150
rect 21170 41620 21210 41660
rect 21830 41650 21870 41690
rect 22070 41650 22110 41690
rect 22310 41650 22350 41690
rect 22550 41650 22590 41690
rect 22790 41650 22830 41690
rect 23030 41650 23070 41690
rect 23270 41650 23310 41690
rect 23510 41650 23550 41690
rect 24430 41760 24470 41800
rect 24670 41760 24710 41800
rect 24910 41760 24950 41800
rect 25150 41760 25190 41800
rect 25390 41760 25430 41800
rect 25630 41760 25670 41800
rect 25870 41760 25910 41800
rect 26110 41760 26150 41800
rect 23950 41540 23990 41580
rect 21160 41270 21200 41310
rect 26280 41270 26320 41310
rect 23950 40920 23990 40960
rect 26270 40870 26320 40920
rect 21160 40610 21200 40650
rect 26480 40620 26520 40660
rect 21160 39520 21200 39560
rect 26730 39520 26770 39560
rect 13210 38920 13250 38960
rect 14210 39040 14260 39090
rect 21830 39060 21870 39100
rect 22070 39060 22110 39100
rect 22310 39060 22350 39100
rect 22550 39060 22590 39100
rect 22790 39060 22830 39100
rect 23030 39060 23070 39100
rect 23270 39060 23310 39100
rect 23510 39060 23550 39100
rect 24430 39170 24470 39210
rect 24670 39170 24710 39210
rect 24910 39170 24950 39210
rect 25150 39170 25190 39210
rect 25390 39170 25430 39210
rect 25630 39170 25670 39210
rect 25870 39170 25910 39210
rect 26110 39170 26150 39210
rect 23950 38950 23990 38990
rect 21160 38830 21200 38870
rect 26480 38840 26520 38880
<< metal1 >>
rect 18430 44100 18530 44110
rect 18430 44020 18440 44100
rect 18520 44020 18530 44100
rect 18430 44010 18530 44020
rect 19170 44100 19270 44110
rect 19170 44020 19180 44100
rect 19260 44020 19270 44100
rect 19170 44010 19270 44020
rect 19910 44100 20010 44110
rect 19910 44020 19920 44100
rect 20000 44020 20010 44100
rect 19910 44010 20010 44020
rect 20650 44100 20750 44110
rect 20650 44020 20660 44100
rect 20740 44020 20750 44100
rect 20650 44010 20750 44020
rect 21390 44100 21490 44110
rect 21390 44020 21400 44100
rect 21480 44020 21490 44100
rect 21390 44010 21490 44020
rect 22130 44100 22230 44110
rect 22130 44020 22140 44100
rect 22220 44020 22230 44100
rect 22130 44010 22230 44020
rect 22870 44100 22970 44110
rect 22870 44020 22880 44100
rect 22960 44020 22970 44100
rect 22870 44010 22970 44020
rect 23590 44100 23690 44110
rect 23590 44020 23600 44100
rect 23680 44020 23690 44100
rect 23590 44010 23690 44020
rect 24350 44100 24490 44110
rect 24350 44020 24360 44100
rect 24440 44020 24490 44100
rect 24350 44010 24490 44020
rect 25090 44100 25190 44110
rect 25090 44020 25100 44100
rect 25180 44020 25190 44100
rect 25090 44010 25190 44020
rect 25830 44100 25930 44110
rect 25830 44020 25840 44100
rect 25920 44020 25930 44100
rect 25830 44010 25930 44020
rect 26570 44100 26670 44110
rect 26570 44020 26580 44100
rect 26660 44020 26670 44100
rect 26570 44010 26670 44020
rect 27310 44100 27410 44110
rect 27310 44020 27320 44100
rect 27400 44020 27410 44100
rect 27310 44010 27410 44020
rect 28050 44100 28150 44110
rect 28050 44020 28060 44100
rect 28140 44020 28150 44100
rect 28050 44010 28150 44020
rect 28790 44100 28890 44110
rect 28790 44020 28800 44100
rect 28880 44020 28890 44100
rect 28790 44010 28890 44020
rect 29530 44100 29630 44110
rect 29530 44020 29540 44100
rect 29620 44020 29630 44100
rect 29530 44010 29630 44020
rect 18470 43690 18530 44010
rect 18470 42650 18550 43690
rect 19210 43680 19270 44010
rect 19200 42830 19280 43680
rect 19950 43660 20010 44010
rect 19940 42990 20020 43660
rect 20690 43650 20750 44010
rect 21430 43650 21490 44010
rect 22170 43680 22230 44010
rect 20680 43160 20760 43650
rect 21420 43350 21500 43650
rect 22160 43520 22240 43680
rect 22910 43660 22970 44010
rect 23630 43660 23690 44010
rect 22910 43580 23330 43660
rect 22160 43440 23090 43520
rect 21420 43270 22850 43350
rect 20680 43080 22610 43160
rect 19940 42910 22370 42990
rect 19200 42750 22130 42830
rect 18470 42570 21890 42650
rect 20880 42220 21280 42230
rect 20880 42040 20890 42220
rect 21070 42150 21280 42220
rect 21070 42110 21160 42150
rect 21200 42110 21280 42150
rect 21070 42040 21280 42110
rect 20880 42030 21280 42040
rect 20880 41720 21280 41730
rect 20880 41540 20890 41720
rect 21070 41660 21280 41720
rect 21070 41620 21170 41660
rect 21210 41620 21280 41660
rect 21070 41540 21280 41620
rect 20880 41530 21280 41540
rect 21810 41690 21890 42570
rect 21810 41650 21830 41690
rect 21870 41650 21890 41690
rect 20880 41380 21280 41390
rect 20880 41200 20890 41380
rect 21070 41310 21280 41380
rect 21070 41270 21160 41310
rect 21200 41270 21280 41310
rect 21070 41200 21280 41270
rect 20880 41190 21280 41200
rect 20870 40710 21270 40720
rect 20870 40530 20880 40710
rect 21060 40650 21270 40710
rect 21060 40610 21160 40650
rect 21200 40610 21270 40650
rect 21060 40530 21270 40610
rect 20870 40520 21270 40530
rect 20880 39630 21280 39640
rect 20880 39450 20890 39630
rect 21070 39560 21280 39630
rect 21070 39520 21160 39560
rect 21200 39520 21280 39560
rect 21070 39450 21280 39520
rect 20880 39440 21280 39450
rect 13189 39073 13271 39374
rect 14168 39110 14410 39120
rect 14168 39090 14300 39110
rect 13190 38960 13270 39073
rect 14168 39066 14210 39090
rect 14170 39040 14210 39066
rect 14260 39040 14300 39090
rect 14170 39010 14300 39040
rect 14400 39010 14410 39110
rect 21810 39100 21890 41650
rect 21810 39060 21830 39100
rect 21870 39060 21890 39100
rect 21810 39040 21890 39060
rect 22050 41690 22130 42750
rect 22050 41650 22070 41690
rect 22110 41650 22130 41690
rect 22050 39100 22130 41650
rect 22050 39060 22070 39100
rect 22110 39060 22130 39100
rect 22050 39040 22130 39060
rect 22290 41690 22370 42910
rect 22290 41650 22310 41690
rect 22350 41650 22370 41690
rect 22290 39100 22370 41650
rect 22290 39060 22310 39100
rect 22350 39060 22370 39100
rect 22290 39040 22370 39060
rect 22530 41690 22610 43080
rect 22530 41650 22550 41690
rect 22590 41650 22610 41690
rect 22530 39100 22610 41650
rect 22530 39060 22550 39100
rect 22590 39060 22610 39100
rect 22530 39040 22610 39060
rect 22770 41690 22850 43270
rect 22770 41650 22790 41690
rect 22830 41650 22850 41690
rect 22770 39100 22850 41650
rect 22770 39060 22790 39100
rect 22830 39060 22850 39100
rect 22770 39040 22850 39060
rect 23010 41690 23090 43440
rect 23010 41650 23030 41690
rect 23070 41650 23090 41690
rect 23010 39100 23090 41650
rect 23010 39060 23030 39100
rect 23070 39060 23090 39100
rect 23010 39040 23090 39060
rect 23250 41690 23330 43580
rect 23250 41650 23270 41690
rect 23310 41650 23330 41690
rect 23250 39100 23330 41650
rect 23250 39060 23270 39100
rect 23310 39060 23330 39100
rect 23250 39040 23330 39060
rect 23490 43580 23690 43660
rect 23490 41690 23570 43580
rect 23490 41650 23510 41690
rect 23550 41650 23570 41690
rect 23490 39100 23570 41650
rect 24410 41800 24490 44010
rect 25130 43660 25190 44010
rect 25870 43660 25930 44010
rect 26610 43660 26670 44010
rect 27350 43670 27410 44010
rect 24410 41760 24430 41800
rect 24470 41760 24490 41800
rect 23930 41580 24010 41600
rect 23930 41561 23950 41580
rect 23929 41540 23950 41561
rect 23990 41561 24010 41580
rect 23990 41540 24011 41561
rect 23929 41073 24011 41540
rect 23930 40960 24010 41073
rect 23930 40920 23950 40960
rect 23990 40920 24010 40960
rect 23930 40900 24010 40920
rect 24410 39210 24490 41760
rect 24410 39170 24430 39210
rect 24470 39170 24490 39210
rect 24410 39150 24490 39170
rect 24650 43580 25190 43660
rect 24650 41800 24730 43580
rect 25850 43520 25930 43660
rect 24650 41760 24670 41800
rect 24710 41760 24730 41800
rect 24650 39210 24730 41760
rect 24650 39170 24670 39210
rect 24710 39170 24730 39210
rect 24650 39150 24730 39170
rect 24890 43440 25930 43520
rect 24890 41800 24970 43440
rect 26600 43350 26680 43660
rect 24890 41760 24910 41800
rect 24950 41760 24970 41800
rect 24890 39210 24970 41760
rect 24890 39170 24910 39210
rect 24950 39170 24970 39210
rect 24890 39150 24970 39170
rect 25130 43270 26680 43350
rect 25130 41800 25210 43270
rect 27340 43170 27420 43670
rect 28090 43660 28150 44010
rect 25130 41760 25150 41800
rect 25190 41760 25210 41800
rect 25130 39210 25210 41760
rect 25130 39170 25150 39210
rect 25190 39170 25210 39210
rect 25130 39150 25210 39170
rect 25370 43090 27420 43170
rect 25370 41800 25450 43090
rect 28070 42970 28150 43660
rect 25370 41760 25390 41800
rect 25430 41760 25450 41800
rect 25370 39210 25450 41760
rect 25370 39170 25390 39210
rect 25430 39170 25450 39210
rect 25370 39150 25450 39170
rect 25610 42890 28150 42970
rect 28830 43700 28890 44010
rect 29570 43720 29630 44010
rect 25610 41800 25690 42890
rect 28830 42840 28910 43700
rect 25610 41760 25630 41800
rect 25670 41760 25690 41800
rect 25610 39210 25690 41760
rect 25610 39170 25630 39210
rect 25670 39170 25690 39210
rect 25610 39150 25690 39170
rect 25850 42760 28910 42840
rect 25850 41800 25930 42760
rect 29570 42660 29650 43720
rect 25850 41760 25870 41800
rect 25910 41760 25930 41800
rect 25850 39210 25930 41760
rect 25850 39170 25870 39210
rect 25910 39170 25930 39210
rect 25850 39150 25930 39170
rect 26090 42580 29650 42660
rect 26090 41800 26170 42580
rect 26650 42220 27050 42230
rect 26650 42150 26860 42220
rect 26650 42110 26730 42150
rect 26770 42110 26860 42150
rect 26650 42040 26860 42110
rect 27040 42040 27050 42220
rect 26650 42030 27050 42040
rect 26090 41760 26110 41800
rect 26150 41760 26170 41800
rect 26090 39210 26170 41760
rect 26200 41380 26600 41390
rect 26200 41310 26410 41380
rect 26200 41270 26280 41310
rect 26320 41270 26410 41310
rect 26200 41200 26410 41270
rect 26590 41200 26600 41380
rect 26200 41190 26600 41200
rect 26240 40940 26470 40950
rect 26240 40920 26360 40940
rect 26240 40870 26270 40920
rect 26320 40870 26360 40920
rect 26240 40840 26360 40870
rect 26460 40840 26470 40940
rect 26240 40830 26470 40840
rect 26410 40660 26610 40730
rect 26410 40620 26480 40660
rect 26520 40620 26610 40660
rect 26410 40520 26610 40620
rect 26410 40340 26420 40520
rect 26600 40340 26610 40520
rect 26410 40330 26610 40340
rect 26650 39630 27050 39640
rect 26650 39560 26860 39630
rect 26650 39520 26730 39560
rect 26770 39520 26860 39560
rect 26650 39450 26860 39520
rect 27040 39450 27050 39630
rect 26650 39440 27050 39450
rect 26090 39170 26110 39210
rect 26150 39170 26170 39210
rect 26090 39150 26170 39170
rect 23490 39060 23510 39100
rect 23550 39060 23570 39100
rect 23490 39040 23570 39060
rect 14170 39000 14410 39010
rect 23930 38990 24010 39010
rect 23930 38971 23950 38990
rect 13190 38920 13210 38960
rect 13250 38920 13270 38960
rect 23929 38950 23950 38971
rect 23990 38971 24010 38990
rect 23990 38950 24011 38971
rect 13190 38900 13270 38920
rect 20870 38930 21270 38940
rect 20870 38750 20880 38930
rect 21060 38870 21270 38930
rect 21060 38830 21160 38870
rect 21200 38830 21270 38870
rect 21060 38750 21270 38830
rect 20870 38740 21270 38750
rect 13270 38470 14010 38480
rect 13270 38370 13900 38470
rect 14000 38370 14010 38470
rect 13270 38360 14010 38370
rect 23929 37730 24011 38950
rect 26410 38880 26610 38950
rect 26410 38840 26480 38880
rect 26520 38840 26610 38880
rect 26410 38740 26610 38840
rect 26410 38560 26420 38740
rect 26600 38560 26610 38740
rect 26410 38550 26610 38560
rect 23910 37720 24030 37730
rect 23910 37620 23920 37720
rect 24020 37620 24030 37720
rect 23910 37610 24030 37620
<< via1 >>
rect 18440 44020 18520 44100
rect 19180 44020 19260 44100
rect 19920 44020 20000 44100
rect 20660 44020 20740 44100
rect 21400 44020 21480 44100
rect 22140 44020 22220 44100
rect 22880 44020 22960 44100
rect 23600 44020 23680 44100
rect 24360 44020 24440 44100
rect 25100 44020 25180 44100
rect 25840 44020 25920 44100
rect 26580 44020 26660 44100
rect 27320 44020 27400 44100
rect 28060 44020 28140 44100
rect 28800 44020 28880 44100
rect 29540 44020 29620 44100
rect 20890 42040 21070 42220
rect 20890 41540 21070 41720
rect 20890 41200 21070 41380
rect 20880 40530 21060 40710
rect 20890 39450 21070 39630
rect 14300 39010 14400 39110
rect 26860 42040 27040 42220
rect 26410 41200 26590 41380
rect 26360 40840 26460 40940
rect 26420 40340 26600 40520
rect 26860 39450 27040 39630
rect 20880 38750 21060 38930
rect 13900 38370 14000 38470
rect 26420 38560 26600 38740
rect 23920 37620 24020 37720
<< metal2 >>
rect 18430 44100 18530 44110
rect 18430 44020 18440 44100
rect 18520 44020 18530 44100
rect 18430 44010 18530 44020
rect 19170 44100 19270 44110
rect 19170 44020 19180 44100
rect 19260 44020 19270 44100
rect 19170 44010 19270 44020
rect 19910 44100 20010 44110
rect 19910 44020 19920 44100
rect 20000 44020 20010 44100
rect 19910 44010 20010 44020
rect 20650 44100 20750 44110
rect 20650 44020 20660 44100
rect 20740 44020 20750 44100
rect 20650 44010 20750 44020
rect 21390 44100 21490 44110
rect 21390 44020 21400 44100
rect 21480 44020 21490 44100
rect 21390 44010 21490 44020
rect 22130 44100 22230 44110
rect 22130 44020 22140 44100
rect 22220 44020 22230 44100
rect 22130 44010 22230 44020
rect 22870 44100 22970 44110
rect 22870 44020 22880 44100
rect 22960 44020 22970 44100
rect 22870 44010 22970 44020
rect 23590 44100 23690 44110
rect 23590 44020 23600 44100
rect 23680 44020 23690 44100
rect 23590 44010 23690 44020
rect 24350 44100 24450 44110
rect 24350 44020 24360 44100
rect 24440 44020 24450 44100
rect 24350 44010 24450 44020
rect 25090 44100 25190 44110
rect 25090 44020 25100 44100
rect 25180 44020 25190 44100
rect 25090 44010 25190 44020
rect 25830 44100 25930 44110
rect 25830 44020 25840 44100
rect 25920 44020 25930 44100
rect 25830 44010 25930 44020
rect 26570 44100 26670 44110
rect 26570 44020 26580 44100
rect 26660 44020 26670 44100
rect 26570 44010 26670 44020
rect 27310 44100 27410 44110
rect 27310 44020 27320 44100
rect 27400 44020 27410 44100
rect 27310 44010 27410 44020
rect 28050 44100 28150 44110
rect 28050 44020 28060 44100
rect 28140 44020 28150 44100
rect 28050 44010 28150 44020
rect 28790 44100 28890 44110
rect 28790 44020 28800 44100
rect 28880 44020 28890 44100
rect 28790 44010 28890 44020
rect 29530 44100 29630 44110
rect 29530 44020 29540 44100
rect 29620 44020 29630 44100
rect 29530 44010 29630 44020
rect 20680 42220 21080 42230
rect 20680 42040 20690 42220
rect 20870 42040 20890 42220
rect 21070 42040 21080 42220
rect 20680 42030 21080 42040
rect 26850 42220 27250 42230
rect 26850 42040 26860 42220
rect 27040 42040 27060 42220
rect 27240 42040 27250 42220
rect 26850 42030 27250 42040
rect 20680 41720 21080 41730
rect 20680 41540 20690 41720
rect 20870 41540 20890 41720
rect 21070 41540 21080 41720
rect 20680 41530 21080 41540
rect 20680 41380 21080 41390
rect 20680 41200 20690 41380
rect 20870 41200 20890 41380
rect 21070 41200 21080 41380
rect 20680 41190 21080 41200
rect 26400 41380 26800 41390
rect 26400 41200 26410 41380
rect 26590 41200 26610 41380
rect 26790 41200 26800 41380
rect 26400 41190 26800 41200
rect 26350 40940 26590 40950
rect 26350 40840 26360 40940
rect 26460 40840 26480 40940
rect 26580 40840 26590 40940
rect 26350 40830 26590 40840
rect 20670 40710 21070 40720
rect 20670 40530 20680 40710
rect 20860 40530 20880 40710
rect 21060 40530 21070 40710
rect 20670 40520 21070 40530
rect 26410 40520 26610 40530
rect 26410 40340 26420 40520
rect 26600 40340 26610 40520
rect 26410 40320 26610 40340
rect 26410 40140 26420 40320
rect 26600 40140 26610 40320
rect 26410 40130 26610 40140
rect 20680 39630 21080 39640
rect 20680 39450 20690 39630
rect 20870 39450 20890 39630
rect 21070 39450 21080 39630
rect 20680 39440 21080 39450
rect 26850 39630 27250 39640
rect 26850 39450 26860 39630
rect 27040 39450 27060 39630
rect 27240 39450 27250 39630
rect 26850 39440 27250 39450
rect 14290 39110 14530 39120
rect 14290 39010 14300 39110
rect 14400 39010 14420 39110
rect 14520 39010 14530 39110
rect 14290 39000 14530 39010
rect 20670 38930 21070 38940
rect 20670 38750 20680 38930
rect 20860 38750 20880 38930
rect 21060 38750 21070 38930
rect 20670 38740 21070 38750
rect 26410 38740 26610 38750
rect 26410 38560 26420 38740
rect 26600 38560 26610 38740
rect 26410 38540 26610 38560
rect 13890 38470 14130 38480
rect 13890 38370 13900 38470
rect 14000 38370 14020 38470
rect 14120 38370 14130 38470
rect 13890 38360 14130 38370
rect 26410 38360 26420 38540
rect 26600 38360 26610 38540
rect 26410 38350 26610 38360
rect 23910 37720 24150 37730
rect 23910 37620 23920 37720
rect 24020 37620 24040 37720
rect 24140 37620 24150 37720
rect 23910 37610 24150 37620
<< rmetal2 >>
rect 18430 44200 18530 44210
rect 18430 44120 18440 44200
rect 18520 44120 18530 44200
rect 18430 44110 18530 44120
rect 19170 44200 19270 44210
rect 19170 44120 19180 44200
rect 19260 44120 19270 44200
rect 19170 44110 19270 44120
rect 19910 44200 20010 44210
rect 19910 44120 19920 44200
rect 20000 44120 20010 44200
rect 19910 44110 20010 44120
rect 20650 44200 20750 44210
rect 20650 44120 20660 44200
rect 20740 44120 20750 44200
rect 20650 44110 20750 44120
rect 21390 44200 21490 44210
rect 21390 44120 21400 44200
rect 21480 44120 21490 44200
rect 21390 44110 21490 44120
rect 22130 44200 22230 44210
rect 22130 44120 22140 44200
rect 22220 44120 22230 44200
rect 22130 44110 22230 44120
rect 22870 44200 22970 44210
rect 22870 44120 22880 44200
rect 22960 44120 22970 44200
rect 22870 44110 22970 44120
rect 23590 44200 23690 44210
rect 23590 44120 23600 44200
rect 23680 44120 23690 44200
rect 23590 44110 23690 44120
rect 24350 44200 24450 44210
rect 24350 44120 24360 44200
rect 24440 44120 24450 44200
rect 24350 44110 24450 44120
rect 25090 44200 25190 44210
rect 25090 44120 25100 44200
rect 25180 44120 25190 44200
rect 25090 44110 25190 44120
rect 25830 44200 25930 44210
rect 25830 44120 25840 44200
rect 25920 44120 25930 44200
rect 25830 44110 25930 44120
rect 26570 44200 26670 44210
rect 26570 44120 26580 44200
rect 26660 44120 26670 44200
rect 26570 44110 26670 44120
rect 27310 44200 27410 44210
rect 27310 44120 27320 44200
rect 27400 44120 27410 44200
rect 27310 44110 27410 44120
rect 28050 44200 28150 44210
rect 28050 44120 28060 44200
rect 28140 44120 28150 44200
rect 28050 44110 28150 44120
rect 28790 44200 28890 44210
rect 28790 44120 28800 44200
rect 28880 44120 28890 44200
rect 28790 44110 28890 44120
rect 29530 44200 29630 44210
rect 29530 44120 29540 44200
rect 29620 44120 29630 44200
rect 29530 44110 29630 44120
<< via2 >>
rect 18440 44120 18520 44200
rect 19180 44120 19260 44200
rect 19920 44120 20000 44200
rect 20660 44120 20740 44200
rect 21400 44120 21480 44200
rect 22140 44120 22220 44200
rect 22880 44120 22960 44200
rect 23600 44120 23680 44200
rect 24360 44120 24440 44200
rect 25100 44120 25180 44200
rect 25840 44120 25920 44200
rect 26580 44120 26660 44200
rect 27320 44120 27400 44200
rect 28060 44120 28140 44200
rect 28800 44120 28880 44200
rect 29540 44120 29620 44200
rect 20690 42040 20870 42220
rect 27060 42040 27240 42220
rect 20690 41540 20870 41720
rect 20690 41200 20870 41380
rect 26610 41200 26790 41380
rect 26480 40840 26580 40940
rect 20680 40530 20860 40710
rect 26420 40140 26600 40320
rect 20690 39450 20870 39630
rect 27060 39450 27240 39630
rect 14420 39010 14520 39110
rect 20680 38750 20860 38930
rect 14020 38370 14120 38470
rect 26420 38360 26600 38540
rect 24040 37620 24140 37720
<< metal3 >>
rect 18430 44300 18530 44310
rect 18430 44220 18440 44300
rect 18520 44220 18530 44300
rect 18430 44200 18530 44220
rect 18430 44120 18440 44200
rect 18520 44120 18530 44200
rect 18430 44110 18530 44120
rect 19170 44300 19270 44310
rect 19170 44220 19180 44300
rect 19260 44220 19270 44300
rect 19170 44200 19270 44220
rect 19170 44120 19180 44200
rect 19260 44120 19270 44200
rect 19170 44110 19270 44120
rect 19910 44300 20010 44310
rect 19910 44220 19920 44300
rect 20000 44220 20010 44300
rect 19910 44200 20010 44220
rect 19910 44120 19920 44200
rect 20000 44120 20010 44200
rect 19910 44110 20010 44120
rect 20650 44300 20750 44310
rect 20650 44220 20660 44300
rect 20740 44220 20750 44300
rect 20650 44200 20750 44220
rect 20650 44120 20660 44200
rect 20740 44120 20750 44200
rect 20650 44110 20750 44120
rect 21390 44300 21490 44310
rect 21390 44220 21400 44300
rect 21480 44220 21490 44300
rect 21390 44200 21490 44220
rect 21390 44120 21400 44200
rect 21480 44120 21490 44200
rect 21390 44110 21490 44120
rect 22130 44300 22230 44310
rect 22130 44220 22140 44300
rect 22220 44220 22230 44300
rect 22130 44200 22230 44220
rect 22130 44120 22140 44200
rect 22220 44120 22230 44200
rect 22130 44110 22230 44120
rect 22870 44300 22970 44310
rect 22870 44220 22880 44300
rect 22960 44220 22970 44300
rect 22870 44200 22970 44220
rect 22870 44120 22880 44200
rect 22960 44120 22970 44200
rect 22870 44110 22970 44120
rect 23590 44300 23690 44310
rect 23590 44220 23600 44300
rect 23680 44220 23690 44300
rect 23590 44200 23690 44220
rect 23590 44120 23600 44200
rect 23680 44120 23690 44200
rect 23590 44110 23690 44120
rect 24350 44300 24450 44310
rect 24350 44220 24360 44300
rect 24440 44220 24450 44300
rect 24350 44200 24450 44220
rect 24350 44120 24360 44200
rect 24440 44120 24450 44200
rect 24350 44110 24450 44120
rect 25090 44300 25190 44310
rect 25090 44220 25100 44300
rect 25180 44220 25190 44300
rect 25090 44200 25190 44220
rect 25090 44120 25100 44200
rect 25180 44120 25190 44200
rect 25090 44110 25190 44120
rect 25830 44300 25930 44310
rect 25830 44220 25840 44300
rect 25920 44220 25930 44300
rect 25830 44200 25930 44220
rect 25830 44120 25840 44200
rect 25920 44120 25930 44200
rect 25830 44110 25930 44120
rect 26570 44300 26670 44310
rect 26570 44220 26580 44300
rect 26660 44220 26670 44300
rect 26570 44200 26670 44220
rect 26570 44120 26580 44200
rect 26660 44120 26670 44200
rect 26570 44110 26670 44120
rect 27310 44300 27410 44310
rect 27310 44220 27320 44300
rect 27400 44220 27410 44300
rect 27310 44200 27410 44220
rect 27310 44120 27320 44200
rect 27400 44120 27410 44200
rect 27310 44110 27410 44120
rect 28050 44300 28150 44310
rect 28050 44220 28060 44300
rect 28140 44220 28150 44300
rect 28050 44200 28150 44220
rect 28050 44120 28060 44200
rect 28140 44120 28150 44200
rect 28050 44110 28150 44120
rect 28790 44300 28890 44310
rect 28790 44220 28800 44300
rect 28880 44220 28890 44300
rect 28790 44200 28890 44220
rect 28790 44120 28800 44200
rect 28880 44120 28890 44200
rect 28790 44110 28890 44120
rect 29530 44300 29630 44310
rect 29530 44220 29540 44300
rect 29620 44220 29630 44300
rect 29530 44200 29630 44220
rect 29530 44120 29540 44200
rect 29620 44120 29630 44200
rect 29530 44110 29630 44120
rect 20390 42310 27310 42570
rect 9280 42270 27310 42310
rect 9280 42220 20880 42270
rect 9280 42040 20690 42220
rect 20870 42040 20880 42220
rect 9280 42010 20880 42040
rect 27010 42220 27310 42270
rect 27010 42040 27060 42220
rect 27240 42040 27310 42220
rect 9280 41470 9580 42010
rect 20480 41720 20880 41730
rect 20480 41540 20490 41720
rect 20670 41540 20690 41720
rect 20870 41540 20880 41720
rect 20480 41530 20880 41540
rect 8898 41460 20880 41470
rect 8898 41180 8910 41460
rect 9190 41380 20880 41460
rect 27010 41450 27310 42040
rect 26540 41390 27310 41450
rect 9190 41200 20690 41380
rect 20870 41200 20880 41380
rect 9190 41180 20880 41200
rect 8898 41170 20880 41180
rect 26560 41380 27310 41390
rect 26560 41200 26610 41380
rect 26790 41200 27310 41380
rect 19730 39720 20030 41170
rect 26560 41140 27310 41200
rect 26470 40940 26710 40950
rect 26470 40840 26480 40940
rect 26580 40840 26600 40940
rect 26700 40840 26710 40940
rect 26470 40830 26710 40840
rect 20470 40710 20870 40720
rect 20470 40530 20480 40710
rect 20660 40530 20680 40710
rect 20860 40530 20870 40710
rect 20470 40520 20870 40530
rect 26410 40320 26610 40330
rect 26410 40140 26420 40320
rect 26600 40140 26610 40320
rect 26410 40120 26610 40140
rect 26410 39940 26420 40120
rect 26600 39940 26610 40120
rect 26410 39930 26610 39940
rect 19730 39630 20880 39720
rect 19730 39450 20690 39630
rect 20870 39450 20880 39630
rect 19730 39420 20880 39450
rect 27000 39630 27310 41140
rect 27000 39450 27060 39630
rect 27240 39450 27310 39630
rect 27000 39445 27310 39450
rect 27010 39440 27310 39445
rect 14410 39110 14650 39120
rect 14410 39010 14420 39110
rect 14520 39010 14540 39110
rect 14640 39010 14650 39110
rect 14410 39000 14650 39010
rect 20480 38930 20870 38940
rect 20660 38750 20680 38930
rect 20860 38750 20870 38930
rect 20480 38740 20870 38750
rect 26410 38540 26610 38550
rect 14010 38470 14250 38480
rect 14010 38370 14020 38470
rect 14120 38370 14140 38470
rect 14240 38370 14250 38470
rect 14010 38360 14250 38370
rect 26410 38360 26420 38540
rect 26600 38360 26610 38540
rect 26410 38340 26610 38360
rect 26410 38160 26420 38340
rect 26600 38160 26610 38340
rect 26410 38150 26610 38160
rect 24030 37720 24270 37730
rect 24030 37620 24040 37720
rect 24140 37620 24160 37720
rect 24260 37620 24270 37720
rect 24030 37610 24270 37620
<< via3 >>
rect 18440 44220 18520 44300
rect 19180 44220 19260 44300
rect 19920 44220 20000 44300
rect 20660 44220 20740 44300
rect 21400 44220 21480 44300
rect 22140 44220 22220 44300
rect 22880 44220 22960 44300
rect 23600 44220 23680 44300
rect 24360 44220 24440 44300
rect 25100 44220 25180 44300
rect 25840 44220 25920 44300
rect 26580 44220 26660 44300
rect 27320 44220 27400 44300
rect 28060 44220 28140 44300
rect 28800 44220 28880 44300
rect 29540 44220 29620 44300
rect 20490 41540 20670 41720
rect 8910 41180 9190 41460
rect 26600 40840 26700 40940
rect 20480 40530 20660 40710
rect 26420 39940 26600 40120
rect 14540 39010 14640 39110
rect 20480 38750 20660 38930
rect 14140 38370 14240 38470
rect 26420 38160 26600 38340
rect 24160 37620 24260 37720
<< metal4 >>
rect 798 44490 858 45152
rect 1534 44490 1594 45152
rect 2270 44490 2330 45152
rect 3006 44490 3066 45152
rect 3742 44490 3802 45152
rect 4478 44490 4538 45152
rect 5214 44490 5274 45152
rect 5950 44490 6010 45152
rect 6686 44490 6746 45152
rect 7422 44490 7482 45152
rect 8158 44490 8218 45152
rect 8894 44490 8954 45152
rect 9630 44490 9690 45152
rect 10366 44490 10426 45152
rect 11102 44490 11162 45152
rect 11838 44490 11898 45152
rect 12574 44490 12634 45152
rect 13310 44490 13370 45152
rect 14046 44490 14106 45152
rect 14782 44490 14842 45152
rect 15518 44490 15578 45152
rect 16254 44490 16314 45152
rect 16990 44490 17050 45152
rect 17726 44490 17786 45152
rect 798 44430 17790 44490
rect 9920 44152 9980 44430
rect 18462 44310 18522 45152
rect 19198 44310 19258 45152
rect 19934 44310 19994 45152
rect 20670 44310 20730 45152
rect 21406 44310 21466 45152
rect 22142 44310 22202 45152
rect 22878 44310 22938 45152
rect 23614 44310 23674 45152
rect 24350 44310 24410 45152
rect 25086 44360 25146 45152
rect 25822 44360 25882 45152
rect 26558 44360 26618 45152
rect 27294 44360 27354 45152
rect 28030 44360 28090 45152
rect 28766 44360 28826 45152
rect 29502 44360 29562 45152
rect 30238 44952 30298 45152
rect 30974 44952 31034 45152
rect 31710 44952 31770 45152
rect 25086 44310 25150 44360
rect 25822 44320 25890 44360
rect 26558 44320 26630 44360
rect 25830 44310 25890 44320
rect 26570 44310 26630 44320
rect 27294 44310 27370 44360
rect 28030 44310 28110 44360
rect 28766 44310 28850 44360
rect 29502 44310 29590 44360
rect 18430 44300 18530 44310
rect 18430 44220 18440 44300
rect 18520 44220 18530 44300
rect 18430 44210 18530 44220
rect 19170 44300 19270 44310
rect 19170 44220 19180 44300
rect 19260 44220 19270 44300
rect 19170 44210 19270 44220
rect 19910 44300 20010 44310
rect 19910 44220 19920 44300
rect 20000 44220 20010 44300
rect 19910 44210 20010 44220
rect 20650 44300 20750 44310
rect 20650 44220 20660 44300
rect 20740 44220 20750 44300
rect 20650 44210 20750 44220
rect 21390 44300 21490 44310
rect 21390 44220 21400 44300
rect 21480 44220 21490 44300
rect 21390 44210 21490 44220
rect 22130 44300 22230 44310
rect 22130 44220 22140 44300
rect 22220 44220 22230 44300
rect 22130 44210 22230 44220
rect 22870 44300 22970 44310
rect 22870 44220 22880 44300
rect 22960 44220 22970 44300
rect 22870 44210 22970 44220
rect 23590 44300 23690 44310
rect 23590 44220 23600 44300
rect 23680 44220 23690 44300
rect 23590 44210 23690 44220
rect 24350 44300 24450 44310
rect 24350 44220 24360 44300
rect 24440 44220 24450 44300
rect 24350 44210 24450 44220
rect 25090 44300 25190 44310
rect 25090 44220 25100 44300
rect 25180 44220 25190 44300
rect 25090 44210 25190 44220
rect 25830 44300 25930 44310
rect 25830 44220 25840 44300
rect 25920 44220 25930 44300
rect 25830 44210 25930 44220
rect 26570 44300 26670 44310
rect 26570 44220 26580 44300
rect 26660 44220 26670 44300
rect 27294 44300 27410 44310
rect 27294 44270 27320 44300
rect 26570 44210 26670 44220
rect 27310 44220 27320 44270
rect 27400 44220 27410 44300
rect 28030 44300 28150 44310
rect 28030 44280 28060 44300
rect 27310 44210 27410 44220
rect 28050 44220 28060 44280
rect 28140 44220 28150 44300
rect 28766 44300 28890 44310
rect 28766 44230 28800 44300
rect 28050 44210 28150 44220
rect 28790 44220 28800 44230
rect 28880 44220 28890 44300
rect 29502 44300 29630 44310
rect 29502 44230 29540 44300
rect 28790 44210 28890 44220
rect 29530 44220 29540 44230
rect 29620 44220 29630 44300
rect 29530 44210 29630 44220
rect 200 41470 500 44152
rect 9800 41808 10100 44152
rect 9800 41720 20680 41808
rect 9800 41540 20490 41720
rect 20670 41540 20680 41720
rect 9800 41508 20680 41540
rect 200 41460 9198 41470
rect 200 41180 8910 41460
rect 9190 41180 9198 41460
rect 200 41170 9198 41180
rect 200 1000 500 41170
rect 9800 40798 10100 41508
rect 26590 40942 26720 40950
rect 26590 40940 31426 40942
rect 26590 40840 26600 40940
rect 26700 40840 31426 40940
rect 26590 40834 31426 40840
rect 26590 40830 26720 40834
rect 9800 40710 20670 40798
rect 9800 40530 20480 40710
rect 20660 40530 20670 40710
rect 9800 40498 20670 40530
rect 9800 1000 10100 40498
rect 20180 40140 20480 40498
rect 20180 40130 26630 40140
rect 20180 40120 26632 40130
rect 20180 39940 26420 40120
rect 26600 39940 26632 40120
rect 20180 39840 26632 39940
rect 14530 39112 14660 39120
rect 14530 39110 14834 39112
rect 14530 39010 14540 39110
rect 14640 39010 14834 39110
rect 14530 39004 14834 39010
rect 20180 39018 20480 39840
rect 14530 39000 14660 39004
rect 20180 38930 20670 39018
rect 20180 38750 20480 38930
rect 20660 38750 20670 38930
rect 20180 38718 20670 38750
rect 14130 38470 14550 38480
rect 14130 38370 14140 38470
rect 14240 38468 14550 38470
rect 14240 38370 14834 38468
rect 14130 38360 14834 38370
rect 14548 38348 14834 38360
rect 20180 38360 20480 38718
rect 20180 38350 26630 38360
rect 20180 38340 26632 38350
rect 20180 38160 26420 38340
rect 26600 38160 26632 38340
rect 20180 38060 26632 38160
rect 24150 37720 27020 37730
rect 24150 37620 24160 37720
rect 24260 37620 27020 37720
rect 24150 37610 27020 37620
rect 26900 34750 27020 37610
rect 26896 34340 27020 34750
rect 400 0 520 200
rect 4816 0 4936 200
rect 9232 0 9352 200
rect 13648 0 13768 200
rect 18064 0 18184 200
rect 22480 0 22600 200
rect 26896 0 27016 34340
rect 31318 34278 31426 40834
rect 31319 200 31425 34278
rect 31312 0 31432 200
<< labels >>
flabel metal4 s 30974 44952 31034 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 31710 44952 31770 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 30238 44952 30298 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 31312 0 31432 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26896 0 27016 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22480 0 22600 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18064 0 18184 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 13648 0 13768 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 9232 0 9352 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 4816 0 4936 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 400 0 520 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 29502 44952 29562 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 28030 44952 28090 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 27294 44952 27354 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 25822 44952 25882 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 25086 44952 25146 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23614 44952 23674 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22878 44952 22938 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21406 44952 21466 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 20670 44952 20730 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19198 44952 19258 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 18462 44952 18522 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 5950 44952 6010 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 5214 44952 5274 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 4478 44952 4538 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 3742 44952 3802 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 3006 44952 3066 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 2270 44952 2330 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 1534 44952 1594 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 798 44952 858 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 10366 44952 10426 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 9630 44952 9690 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 8158 44952 8218 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 7422 44952 7482 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 16990 44952 17050 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 16254 44952 16314 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 14782 44952 14842 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 14046 44952 14106 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 12574 44952 12634 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 11838 44952 11898 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 200 1000 500 44152 1 FreeSans 2 0 0 0 VPWR
port 51 nsew power bidirectional
rlabel viali 23950 41540 23990 41580 1 Idiff
flabel metal4 9800 1000 10100 44152 1 FreeSans 2 0 0 0 VGND
port 52 nsew ground bidirectional
rlabel viali 23950 38950 23990 38990 1 Idiff
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
