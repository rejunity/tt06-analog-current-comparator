Current Comparator Simulation
* this file edited to remove everything not in tt lib
* .lib "./sky130_fd_pr/models/sky130.lib.spice" tt
.lib "/Users/rej/.volare/sky130A/libs.tech/ngspice/sky130.lib.spice" tt

* instantiate the Current Comparator
Xinv Y A VGND VPWR tt_um_rejunity_current_cmp

.subckt tt_um_rejunity_current_cmp Y A VGND VPWR
* NGSPICE file created from tt_um_rejunity_current_cmp.ext - technology: sky130A

X0 Y A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.189 pd=1.74 as=0.168 ps=1.64 w=0.42 l=0.15
X1 Y A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.45 pd=2.9 as=0.4 ps=2.8 w=1 l=0.15
C15 m3_201_22427# VPWR 0.40909f
C16 Y VPWR 0.098215f
C18 A VPWR 0.048717f
C20 A Y 0.036438f
C113 VPWR VGND 24.929401f
C114 m3_201_22427# VGND 4.47465f $ **FLOATING
C115 Y VGND 0.185356f
C116 A VGND 0.301948f


.ends

* set gnd and power
Vgnd VGND 0 0
Vdd VPWR VGND 1.8

* create pulse
Vin A VGND pulse(0 1.8 1p 10p 10p 1n 2n)
.tran 10e-12 2e-09 0e-00

.control
run
set color0 = white
set color1 = black
plot A Y
plot i(Vdd)
.endc

.end
