* NGSPICE file created from tt_um_rejunity_current_cmp.ext - technology: sky130A

.subckt tt_um_rejunity_current_cmp clk ena rst_n ua[0] ua[1] ua[2] ua[3] ua[4] ua[5]
+ ua[6] ua[7] ui_in[0] ui_in[1] ui_in[2] ui_in[3] ui_in[4] ui_in[5] ui_in[6] ui_in[7]
+ uio_in[0] uio_in[1] uio_in[2] uio_in[3] uio_in[4] uio_in[5] uio_in[6] uio_in[7]
+ uio_oe[0] uio_oe[1] uio_oe[2] uio_oe[3] uio_oe[4] uio_oe[5] uio_oe[6] uio_oe[7]
+ uio_out[0] uio_out[1] uio_out[2] uio_out[3] uio_out[4] uio_out[5] uio_out[6] uio_out[7]
+ uo_out[0] uo_out[1] uo_out[2] uo_out[3] uo_out[4] uo_out[5] uo_out[6] uo_out[7]
+ VPWR VGND
X0 Y A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.189 pd=1.74 as=0.168 ps=1.64 w=0.42 l=0.15
**devattr s=6720,328 d=7560,348
X1 Y A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.45 pd=2.9 as=0.4 ps=2.8 w=1 l=0.15
**devattr s=16000,560 d=18000,580
.ends

