magic
tech sky130A
magscale 1 2
timestamp 1713440464
<< nwell >>
rect 12360 43810 14180 44190
rect 12870 42970 13600 43350
<< nmos >>
rect 12580 43520 12610 43604
rect 12820 43520 12850 43604
rect 13460 43520 13490 43604
rect 13740 43520 13770 43604
rect 13980 43520 14010 43604
rect 13070 42710 13100 42794
rect 13400 42710 13430 42794
<< pmos >>
rect 12580 43850 12610 44050
rect 12820 43850 12850 44050
rect 13140 43850 13170 44050
rect 13740 43850 13770 44050
rect 13980 43850 14010 44050
rect 13070 43010 13100 43210
rect 13400 43010 13430 43210
<< ndiff >>
rect 12500 43580 12580 43604
rect 12500 43540 12520 43580
rect 12560 43540 12580 43580
rect 12500 43520 12580 43540
rect 12610 43580 12680 43604
rect 12610 43540 12630 43580
rect 12670 43540 12680 43580
rect 12610 43520 12680 43540
rect 12740 43580 12820 43604
rect 12740 43540 12760 43580
rect 12800 43540 12820 43580
rect 12740 43520 12820 43540
rect 12850 43580 12920 43604
rect 12850 43540 12870 43580
rect 12910 43540 12920 43580
rect 12850 43520 12920 43540
rect 13350 43580 13460 43604
rect 13350 43540 13360 43580
rect 13440 43540 13460 43580
rect 13350 43520 13460 43540
rect 13490 43580 13600 43604
rect 13490 43540 13510 43580
rect 13590 43540 13600 43580
rect 13490 43520 13600 43540
rect 13660 43580 13740 43604
rect 13660 43540 13680 43580
rect 13720 43540 13740 43580
rect 13660 43520 13740 43540
rect 13770 43580 13840 43604
rect 13770 43540 13790 43580
rect 13830 43540 13840 43580
rect 13770 43520 13840 43540
rect 13900 43580 13980 43604
rect 13900 43540 13920 43580
rect 13960 43540 13980 43580
rect 13900 43520 13980 43540
rect 14010 43580 14080 43604
rect 14010 43540 14030 43580
rect 14070 43540 14080 43580
rect 14010 43520 14080 43540
rect 12980 42770 13070 42794
rect 12980 42730 13010 42770
rect 13050 42730 13070 42770
rect 12980 42710 13070 42730
rect 13100 42770 13180 42794
rect 13100 42730 13120 42770
rect 13160 42730 13180 42770
rect 13100 42710 13180 42730
rect 13320 42770 13400 42794
rect 13320 42730 13340 42770
rect 13380 42730 13400 42770
rect 13320 42710 13400 42730
rect 13430 42770 13520 42794
rect 13430 42730 13450 42770
rect 13490 42730 13520 42770
rect 13430 42710 13520 42730
<< pdiff >>
rect 12500 44020 12580 44050
rect 12500 43880 12520 44020
rect 12560 43880 12580 44020
rect 12500 43850 12580 43880
rect 12610 44020 12680 44050
rect 12610 43880 12630 44020
rect 12670 43880 12680 44020
rect 12610 43850 12680 43880
rect 12740 44020 12820 44050
rect 12740 43880 12760 44020
rect 12800 43880 12820 44020
rect 12740 43850 12820 43880
rect 12850 44020 12920 44050
rect 12850 43880 12870 44020
rect 12910 43880 12920 44020
rect 12850 43850 12920 43880
rect 13030 44020 13140 44050
rect 13030 43880 13040 44020
rect 13120 43880 13140 44020
rect 13030 43850 13140 43880
rect 13170 44020 13280 44050
rect 13170 43880 13190 44020
rect 13270 43880 13280 44020
rect 13170 43850 13280 43880
rect 13660 44020 13740 44050
rect 13660 43880 13680 44020
rect 13720 43880 13740 44020
rect 13660 43850 13740 43880
rect 13770 44020 13840 44050
rect 13770 43880 13790 44020
rect 13830 43880 13840 44020
rect 13770 43850 13840 43880
rect 13900 44020 13980 44050
rect 13900 43880 13920 44020
rect 13960 43880 13980 44020
rect 13900 43850 13980 43880
rect 14010 44020 14080 44050
rect 14010 43880 14030 44020
rect 14070 43880 14080 44020
rect 14010 43850 14080 43880
rect 12910 43180 13070 43210
rect 12910 43040 12930 43180
rect 12970 43040 13070 43180
rect 12910 43010 13070 43040
rect 13100 43180 13180 43210
rect 13100 43040 13120 43180
rect 13160 43040 13180 43180
rect 13100 43010 13180 43040
rect 13320 43180 13400 43210
rect 13320 43040 13340 43180
rect 13380 43040 13400 43180
rect 13320 43010 13400 43040
rect 13430 43180 13520 43210
rect 13430 43040 13450 43180
rect 13490 43040 13520 43180
rect 13430 43010 13520 43040
<< ndiffc >>
rect 12520 43540 12560 43580
rect 12630 43540 12670 43580
rect 12760 43540 12800 43580
rect 12870 43540 12910 43580
rect 13360 43540 13440 43580
rect 13510 43540 13590 43580
rect 13680 43540 13720 43580
rect 13790 43540 13830 43580
rect 13920 43540 13960 43580
rect 14030 43540 14070 43580
rect 13010 42730 13050 42770
rect 13120 42730 13160 42770
rect 13340 42730 13380 42770
rect 13450 42730 13490 42770
<< pdiffc >>
rect 12520 43880 12560 44020
rect 12630 43880 12670 44020
rect 12760 43880 12800 44020
rect 12870 43880 12910 44020
rect 13040 43880 13120 44020
rect 13190 43880 13270 44020
rect 13680 43880 13720 44020
rect 13790 43880 13830 44020
rect 13920 43880 13960 44020
rect 14030 43880 14070 44020
rect 12930 43040 12970 43180
rect 13120 43040 13160 43180
rect 13340 43040 13380 43180
rect 13450 43040 13490 43180
<< psubdiff >>
rect 12400 43420 12430 43460
rect 12470 43420 12500 43460
rect 12560 43420 12590 43460
rect 12630 43420 12660 43460
rect 12720 43420 12750 43460
rect 12790 43420 12820 43460
rect 12880 43420 12910 43460
rect 12950 43420 12980 43460
rect 13400 43420 13430 43460
rect 13470 43420 13500 43460
rect 13560 43420 13590 43460
rect 13630 43420 13660 43460
rect 13720 43420 13750 43460
rect 13790 43420 13820 43460
rect 13880 43420 13910 43460
rect 13950 43420 13980 43460
rect 14040 43420 14070 43460
rect 14110 43420 14140 43460
rect 12980 42610 13010 42650
rect 13050 42610 13080 42650
rect 13140 42610 13170 42650
rect 13210 42610 13240 42650
rect 13300 42610 13330 42650
rect 13370 42610 13400 42650
rect 13460 42610 13490 42650
rect 13530 42610 13560 42650
<< nsubdiff >>
rect 12400 44110 12430 44150
rect 12470 44110 12500 44150
rect 12560 44110 12590 44150
rect 12630 44110 12660 44150
rect 12720 44110 12750 44150
rect 12790 44110 12820 44150
rect 12880 44110 12910 44150
rect 12950 44110 12980 44150
rect 13040 44110 13070 44150
rect 13110 44110 13140 44150
rect 13200 44110 13230 44150
rect 13270 44110 13300 44150
rect 13560 44110 13590 44150
rect 13630 44110 13660 44150
rect 13720 44110 13750 44150
rect 13790 44110 13820 44150
rect 13880 44110 13910 44150
rect 13950 44110 13980 44150
rect 14040 44110 14070 44150
rect 14110 44110 14140 44150
rect 12980 43270 13010 43310
rect 13050 43270 13080 43310
rect 13140 43270 13170 43310
rect 13210 43270 13240 43310
rect 13300 43270 13330 43310
rect 13370 43270 13400 43310
rect 13460 43270 13490 43310
rect 13530 43270 13560 43310
<< psubdiffcont >>
rect 12430 43420 12470 43460
rect 12590 43420 12630 43460
rect 12750 43420 12790 43460
rect 12910 43420 12950 43460
rect 13430 43420 13470 43460
rect 13590 43420 13630 43460
rect 13750 43420 13790 43460
rect 13910 43420 13950 43460
rect 14070 43420 14110 43460
rect 13010 42610 13050 42650
rect 13170 42610 13210 42650
rect 13330 42610 13370 42650
rect 13490 42610 13530 42650
<< nsubdiffcont >>
rect 12430 44110 12470 44150
rect 12590 44110 12630 44150
rect 12750 44110 12790 44150
rect 12910 44110 12950 44150
rect 13070 44110 13110 44150
rect 13230 44110 13270 44150
rect 13590 44110 13630 44150
rect 13750 44110 13790 44150
rect 13910 44110 13950 44150
rect 14070 44110 14110 44150
rect 13010 43270 13050 43310
rect 13170 43270 13210 43310
rect 13330 43270 13370 43310
rect 13490 43270 13530 43310
<< poly >>
rect 12580 44050 12610 44080
rect 12820 44050 12850 44080
rect 13140 44050 13170 44080
rect 13740 44050 13770 44080
rect 13980 44050 14010 44080
rect 12580 43810 12610 43850
rect 12820 43810 12850 43850
rect 13140 43810 13170 43850
rect 13740 43810 13770 43850
rect 13980 43810 14010 43850
rect 12580 43800 12690 43810
rect 12580 43760 12630 43800
rect 12670 43760 12690 43800
rect 12580 43750 12690 43760
rect 12820 43800 12930 43810
rect 12820 43760 12870 43800
rect 12910 43760 12930 43800
rect 12820 43750 12930 43760
rect 13030 43800 13170 43810
rect 13030 43720 13050 43800
rect 13130 43720 13170 43800
rect 13670 43800 13770 43810
rect 13670 43760 13690 43800
rect 13730 43760 13770 43800
rect 13670 43750 13770 43760
rect 13910 43800 14010 43810
rect 13910 43760 13930 43800
rect 13970 43760 14010 43800
rect 13910 43750 14010 43760
rect 13030 43710 13170 43720
rect 13460 43720 13590 43730
rect 12510 43690 12610 43700
rect 12510 43650 12530 43690
rect 12570 43650 12610 43690
rect 12510 43640 12610 43650
rect 12750 43690 12850 43700
rect 12750 43650 12770 43690
rect 12810 43650 12850 43690
rect 12750 43640 12850 43650
rect 12580 43604 12610 43640
rect 12820 43604 12850 43640
rect 13460 43650 13500 43720
rect 13570 43650 13590 43720
rect 13460 43640 13590 43650
rect 13740 43690 13830 43700
rect 13740 43650 13770 43690
rect 13810 43650 13830 43690
rect 13740 43640 13830 43650
rect 13980 43690 14070 43700
rect 13980 43650 14010 43690
rect 14050 43650 14070 43690
rect 13980 43640 14070 43650
rect 13460 43604 13490 43640
rect 13740 43604 13770 43640
rect 13980 43604 14010 43640
rect 12580 43490 12610 43520
rect 12820 43490 12850 43520
rect 13460 43490 13490 43520
rect 13740 43490 13770 43520
rect 13980 43490 14010 43520
rect 13070 43210 13100 43240
rect 13400 43210 13430 43240
rect 13070 42890 13100 43010
rect 13400 42970 13430 43010
rect 13320 42960 13430 42970
rect 13320 42920 13340 42960
rect 13380 42920 13430 42960
rect 13320 42910 13430 42920
rect 13070 42880 13280 42890
rect 13070 42840 13220 42880
rect 13260 42840 13280 42880
rect 13070 42830 13280 42840
rect 13070 42794 13100 42830
rect 13400 42794 13430 42910
rect 13070 42680 13100 42710
rect 13400 42680 13430 42710
<< polycont >>
rect 12630 43760 12670 43800
rect 12870 43760 12910 43800
rect 13050 43720 13130 43800
rect 13690 43760 13730 43800
rect 13930 43760 13970 43800
rect 12530 43650 12570 43690
rect 12770 43650 12810 43690
rect 13500 43650 13570 43720
rect 13770 43650 13810 43690
rect 14010 43650 14050 43690
rect 13340 42920 13380 42960
rect 13220 42840 13260 42880
<< locali >>
rect 11530 44150 14150 44170
rect 11530 44110 12430 44150
rect 12470 44110 12590 44150
rect 12630 44110 12750 44150
rect 12790 44110 12910 44150
rect 12950 44110 13070 44150
rect 13110 44110 13230 44150
rect 13270 44110 13590 44150
rect 13630 44110 13750 44150
rect 13790 44110 13910 44150
rect 13950 44110 14070 44150
rect 14110 44110 14150 44150
rect 11530 44090 14150 44110
rect 11530 43990 11610 44090
rect 11000 43970 11610 43990
rect 11000 43930 11020 43970
rect 11060 43930 11610 43970
rect 11000 43910 11610 43930
rect 12500 44020 12560 44090
rect 12500 43880 12520 44020
rect 12500 43850 12560 43880
rect 12630 44020 12670 44050
rect 12630 43810 12670 43880
rect 12740 44020 12800 44090
rect 12740 43880 12760 44020
rect 12740 43850 12800 43880
rect 12870 44020 12910 44050
rect 12870 43810 12910 43880
rect 13040 44020 13120 44090
rect 13040 43850 13120 43880
rect 13190 44020 13270 44050
rect 12440 43800 13150 43810
rect 12440 43760 12630 43800
rect 12670 43760 12870 43800
rect 12910 43760 13050 43800
rect 12440 43730 13050 43760
rect 11010 43660 11610 43680
rect 11010 43620 11030 43660
rect 11070 43620 11610 43660
rect 12510 43650 12530 43690
rect 12570 43650 12590 43690
rect 11010 43600 11610 43620
rect 11530 43480 11610 43600
rect 12500 43580 12560 43600
rect 12500 43540 12520 43580
rect 12500 43480 12560 43540
rect 12630 43580 12670 43730
rect 12870 43720 13050 43730
rect 13130 43720 13150 43800
rect 12870 43710 13150 43720
rect 12750 43650 12770 43690
rect 12810 43650 12830 43690
rect 12630 43520 12670 43540
rect 12740 43580 12800 43600
rect 12740 43540 12760 43580
rect 12740 43480 12800 43540
rect 12870 43580 12910 43710
rect 12870 43520 12910 43540
rect 13190 43600 13270 43880
rect 13660 44020 13720 44090
rect 13660 43880 13680 44020
rect 13660 43850 13720 43880
rect 13790 44020 13830 44050
rect 13670 43800 13750 43810
rect 13670 43760 13690 43800
rect 13730 43760 13750 43800
rect 13670 43750 13750 43760
rect 13480 43720 13590 43730
rect 13480 43650 13500 43720
rect 13570 43710 13590 43720
rect 13790 43710 13830 43880
rect 13900 44020 13960 44090
rect 13900 43880 13920 44020
rect 13900 43850 13960 43880
rect 14030 44020 14070 44050
rect 13910 43800 13990 43810
rect 13910 43760 13930 43800
rect 13970 43760 13990 43800
rect 13910 43750 13990 43760
rect 14030 43710 14070 43880
rect 13570 43690 14070 43710
rect 13570 43650 13770 43690
rect 13810 43650 14010 43690
rect 14050 43650 14070 43690
rect 13480 43640 14070 43650
rect 13190 43580 13440 43600
rect 13190 43540 13210 43580
rect 13250 43540 13360 43580
rect 13190 43520 13440 43540
rect 13510 43580 13590 43600
rect 13510 43480 13590 43540
rect 13680 43580 13720 43600
rect 13680 43480 13720 43540
rect 13790 43580 13830 43640
rect 13790 43520 13830 43540
rect 13900 43580 13960 43600
rect 13900 43540 13920 43580
rect 13900 43480 13960 43540
rect 14030 43580 14070 43640
rect 14030 43520 14070 43540
rect 11530 43460 14130 43480
rect 11530 43420 12430 43460
rect 12470 43420 12590 43460
rect 12630 43420 12750 43460
rect 12790 43420 12910 43460
rect 12950 43420 13430 43460
rect 13470 43420 13590 43460
rect 13630 43420 13750 43460
rect 13790 43420 13910 43460
rect 13950 43420 14070 43460
rect 14110 43420 14130 43460
rect 11530 43400 14130 43420
rect 11000 43310 13550 43330
rect 11000 43270 11020 43310
rect 11060 43270 13010 43310
rect 13050 43270 13170 43310
rect 13210 43270 13330 43310
rect 13370 43270 13490 43310
rect 13530 43270 13550 43310
rect 11000 43250 13550 43270
rect 12930 43180 12970 43210
rect 12930 42670 12970 43040
rect 13010 42770 13050 43250
rect 13010 42710 13050 42730
rect 13120 43180 13160 43210
rect 13120 42960 13160 43040
rect 13320 43180 13380 43250
rect 13320 43040 13340 43180
rect 13320 43010 13380 43040
rect 13450 43180 13510 43210
rect 13490 43040 13510 43180
rect 13120 42920 13210 42960
rect 13250 42920 13340 42960
rect 13380 42920 13400 42960
rect 13450 42920 13510 43040
rect 13810 42920 13860 43040
rect 13120 42770 13160 42920
rect 13450 42880 13860 42920
rect 13200 42840 13220 42880
rect 13260 42840 13510 42880
rect 13120 42710 13160 42730
rect 13320 42770 13380 42790
rect 13320 42730 13340 42770
rect 13320 42670 13380 42730
rect 13450 42770 13510 42840
rect 13490 42730 13510 42770
rect 13450 42710 13510 42730
rect 11010 42650 13550 42670
rect 11010 42610 11030 42650
rect 11070 42610 13010 42650
rect 13050 42610 13170 42650
rect 13210 42610 13330 42650
rect 13370 42610 13490 42650
rect 13530 42610 13550 42650
rect 11010 42590 13550 42610
<< viali >>
rect 11020 43930 11060 43970
rect 11030 43620 11070 43660
rect 12530 43650 12570 43690
rect 12770 43650 12810 43690
rect 13690 43760 13730 43800
rect 13930 43760 13970 43800
rect 13210 43540 13250 43580
rect 11020 43270 11060 43310
rect 13210 42920 13250 42960
rect 13810 43040 13860 43090
rect 11030 42610 11070 42650
<< metal1 >>
rect 22140 44460 22240 44470
rect 22140 44430 22150 44460
rect 12510 44380 22150 44430
rect 22230 44380 22240 44460
rect 12510 44370 22240 44380
rect 22460 44370 22560 44380
rect 10740 44040 11140 44050
rect 10740 43860 10750 44040
rect 10930 43970 11140 44040
rect 10930 43930 11020 43970
rect 11060 43930 11140 43970
rect 10930 43860 11140 43930
rect 10740 43850 11140 43860
rect 10740 43720 11140 43730
rect 10740 43540 10750 43720
rect 10930 43660 11140 43720
rect 10930 43620 11030 43660
rect 11070 43620 11140 43660
rect 12510 43690 12590 44370
rect 22460 44340 22470 44370
rect 12510 43650 12530 43690
rect 12570 43650 12590 43690
rect 12510 43630 12590 43650
rect 12750 44290 22470 44340
rect 22550 44290 22560 44370
rect 12750 44280 22560 44290
rect 23740 44280 23840 44290
rect 12750 43690 12830 44280
rect 23740 44250 23750 44280
rect 13670 44200 23750 44250
rect 23830 44200 23840 44280
rect 13670 44190 23840 44200
rect 24060 44190 24160 44200
rect 13670 43800 13750 44190
rect 24060 44160 24070 44190
rect 14230 44110 24070 44160
rect 24150 44110 24160 44190
rect 14230 44100 24160 44110
rect 14230 43820 14310 44100
rect 13670 43760 13690 43800
rect 13730 43760 13750 43800
rect 13670 43740 13750 43760
rect 13910 43800 14310 43820
rect 13910 43760 13930 43800
rect 13970 43760 14310 43800
rect 13910 43740 14310 43760
rect 12750 43650 12770 43690
rect 12810 43650 12830 43690
rect 12750 43630 12830 43650
rect 10930 43540 11140 43620
rect 10740 43530 11140 43540
rect 13190 43580 13270 43600
rect 13190 43540 13210 43580
rect 13250 43540 13270 43580
rect 10740 43380 11140 43390
rect 10740 43200 10750 43380
rect 10930 43310 11140 43380
rect 10930 43270 11020 43310
rect 11060 43270 11140 43310
rect 10930 43200 11140 43270
rect 10740 43190 11140 43200
rect 13190 42960 13270 43540
rect 13770 43110 14010 43120
rect 13770 43090 13900 43110
rect 13770 43040 13810 43090
rect 13860 43040 13900 43090
rect 13770 43010 13900 43040
rect 14000 43010 14010 43110
rect 13770 43000 14010 43010
rect 13190 42920 13210 42960
rect 13250 42920 13270 42960
rect 13190 42900 13270 42920
rect 10740 42710 11140 42720
rect 10740 42530 10750 42710
rect 10930 42650 11140 42710
rect 10930 42610 11030 42650
rect 11070 42610 11140 42650
rect 10930 42530 11140 42610
rect 10740 42520 11140 42530
rect 13270 42470 14010 42480
rect 13270 42370 13900 42470
rect 14000 42370 14010 42470
rect 13270 42360 14010 42370
<< via1 >>
rect 22150 44380 22230 44460
rect 10750 43860 10930 44040
rect 10750 43540 10930 43720
rect 22470 44290 22550 44370
rect 23750 44200 23830 44280
rect 24070 44110 24150 44190
rect 10750 43200 10930 43380
rect 13900 43010 14000 43110
rect 10750 42530 10930 42710
rect 13900 42370 14000 42470
<< metal2 >>
rect 22140 44460 22240 44470
rect 22140 44380 22150 44460
rect 22230 44380 22240 44460
rect 22140 44370 22240 44380
rect 22460 44370 22560 44380
rect 22460 44290 22470 44370
rect 22550 44290 22560 44370
rect 22460 44280 22560 44290
rect 23740 44280 23840 44290
rect 23740 44200 23750 44280
rect 23830 44200 23840 44280
rect 23740 44190 23840 44200
rect 24060 44190 24160 44200
rect 24060 44110 24070 44190
rect 24150 44110 24160 44190
rect 24060 44100 24160 44110
rect 10540 44040 10940 44050
rect 10540 43860 10550 44040
rect 10730 43860 10750 44040
rect 10930 43860 10940 44040
rect 10540 43850 10940 43860
rect 10540 43720 10940 43730
rect 10540 43540 10550 43720
rect 10730 43540 10750 43720
rect 10930 43540 10940 43720
rect 10540 43530 10940 43540
rect 10540 43380 10940 43390
rect 10540 43200 10550 43380
rect 10730 43200 10750 43380
rect 10930 43200 10940 43380
rect 10540 43190 10940 43200
rect 13890 43110 14130 43120
rect 13890 43010 13900 43110
rect 14000 43010 14020 43110
rect 14120 43010 14130 43110
rect 13890 43000 14130 43010
rect 10540 42710 10940 42720
rect 10540 42530 10550 42710
rect 10730 42530 10750 42710
rect 10930 42530 10940 42710
rect 10540 42520 10940 42530
rect 13890 42470 14130 42480
rect 13890 42370 13900 42470
rect 14000 42370 14020 42470
rect 14120 42370 14130 42470
rect 13890 42360 14130 42370
<< rmetal2 >>
rect 22240 44460 22340 44470
rect 22240 44380 22250 44460
rect 22330 44380 22340 44460
rect 22240 44370 22340 44380
rect 22560 44370 22660 44380
rect 22560 44290 22570 44370
rect 22650 44290 22660 44370
rect 22560 44280 22660 44290
rect 23840 44280 23940 44290
rect 23840 44200 23850 44280
rect 23930 44200 23940 44280
rect 23840 44190 23940 44200
rect 24160 44190 24260 44200
rect 24160 44110 24170 44190
rect 24250 44110 24260 44190
rect 24160 44100 24260 44110
<< via2 >>
rect 22250 44380 22330 44460
rect 22570 44290 22650 44370
rect 23850 44200 23930 44280
rect 24170 44110 24250 44190
rect 10550 43860 10730 44040
rect 10550 43540 10730 43720
rect 10550 43200 10730 43380
rect 14020 43010 14120 43110
rect 10550 42530 10730 42710
rect 14020 42370 14120 42470
<< metal3 >>
rect 22240 44460 22440 44470
rect 22240 44380 22250 44460
rect 22330 44380 22350 44460
rect 22430 44380 22440 44460
rect 22240 44370 22440 44380
rect 22560 44370 22760 44380
rect 22560 44290 22570 44370
rect 22650 44290 22670 44370
rect 22750 44290 22760 44370
rect 22560 44280 22760 44290
rect 23840 44280 24040 44290
rect 23840 44200 23850 44280
rect 23930 44200 23950 44280
rect 24030 44200 24040 44280
rect 23840 44190 24040 44200
rect 24160 44190 24360 44200
rect 9280 44040 10740 44130
rect 24160 44110 24170 44190
rect 24250 44110 24270 44190
rect 24350 44110 24360 44190
rect 24160 44100 24360 44110
rect 9280 43860 10550 44040
rect 10730 43860 10740 44040
rect 9280 43830 10740 43860
rect 9280 43470 9580 43830
rect 10340 43720 10740 43730
rect 10340 43540 10350 43720
rect 10530 43540 10550 43720
rect 10730 43540 10740 43720
rect 10340 43530 10740 43540
rect 8898 43460 10740 43470
rect 8898 43180 8910 43460
rect 9190 43380 10740 43460
rect 9190 43200 10550 43380
rect 10730 43200 10740 43380
rect 9190 43180 10740 43200
rect 8898 43170 10740 43180
rect 14010 43110 14250 43120
rect 14010 43010 14020 43110
rect 14120 43010 14140 43110
rect 14240 43010 14250 43110
rect 14010 43000 14250 43010
rect 10340 42710 10740 42720
rect 10340 42530 10350 42710
rect 10530 42530 10550 42710
rect 10730 42530 10740 42710
rect 10340 42520 10740 42530
rect 14010 42470 14250 42480
rect 14010 42370 14020 42470
rect 14120 42370 14140 42470
rect 14240 42370 14250 42470
rect 14010 42360 14250 42370
<< via3 >>
rect 22350 44380 22430 44460
rect 22670 44290 22750 44370
rect 23950 44200 24030 44280
rect 24270 44110 24350 44190
rect 10350 43540 10530 43720
rect 8910 43180 9190 43460
rect 14140 43010 14240 43110
rect 10350 42530 10530 42710
rect 14140 42370 14240 42470
<< metal4 >>
rect 798 44490 858 45152
rect 1534 44490 1594 45152
rect 2270 44490 2330 45152
rect 3006 44490 3066 45152
rect 3742 44490 3802 45152
rect 4478 44490 4538 45152
rect 5214 44490 5274 45152
rect 5950 44490 6010 45152
rect 6686 44490 6746 45152
rect 7422 44490 7482 45152
rect 8158 44490 8218 45152
rect 8894 44490 8954 45152
rect 9630 44490 9690 45152
rect 10366 44490 10426 45152
rect 11102 44490 11162 45152
rect 11838 44490 11898 45152
rect 12574 44490 12634 45152
rect 13310 44490 13370 45152
rect 14046 44490 14106 45152
rect 14782 44490 14842 45152
rect 15518 44490 15578 45152
rect 16254 44490 16314 45152
rect 16990 44490 17050 45152
rect 17726 44490 17786 45152
rect 18462 44952 18522 45152
rect 19198 44952 19258 45152
rect 19934 44952 19994 45152
rect 20670 44952 20730 45152
rect 21406 44952 21466 45152
rect 22142 44952 22202 45152
rect 22878 44530 22938 45152
rect 798 44430 17790 44490
rect 22340 44470 22938 44530
rect 22340 44460 22440 44470
rect 9920 44152 9980 44430
rect 22340 44380 22350 44460
rect 22430 44380 22440 44460
rect 23614 44380 23674 45152
rect 22340 44370 22440 44380
rect 22660 44370 23674 44380
rect 22660 44290 22670 44370
rect 22750 44320 23674 44370
rect 24350 44350 24410 45152
rect 22750 44290 22760 44320
rect 22660 44280 22760 44290
rect 23940 44290 24410 44350
rect 23940 44280 24040 44290
rect 23940 44200 23950 44280
rect 24030 44200 24040 44280
rect 25086 44200 25146 45152
rect 25822 44952 25882 45152
rect 26558 44952 26618 45152
rect 27294 44952 27354 45152
rect 28030 44952 28090 45152
rect 28766 44952 28826 45152
rect 29502 44952 29562 45152
rect 30238 44952 30298 45152
rect 30974 44952 31034 45152
rect 31710 44952 31770 45152
rect 23940 44190 24040 44200
rect 24260 44190 25146 44200
rect 200 43470 500 44152
rect 9800 43808 10100 44152
rect 24260 44110 24270 44190
rect 24350 44140 25146 44190
rect 24350 44110 24360 44140
rect 24260 44100 24360 44110
rect 9800 43720 10540 43808
rect 9800 43540 10350 43720
rect 10530 43540 10540 43720
rect 9800 43508 10540 43540
rect 200 43460 9198 43470
rect 200 43180 8910 43460
rect 9190 43180 9198 43460
rect 200 43170 9198 43180
rect 200 1000 500 43170
rect 9800 42798 10100 43508
rect 14130 43112 14260 43120
rect 14130 43110 31426 43112
rect 14130 43010 14140 43110
rect 14240 43010 31426 43110
rect 14130 43004 31426 43010
rect 14130 43000 14260 43004
rect 9800 42710 10540 42798
rect 9800 42530 10350 42710
rect 10530 42530 10540 42710
rect 9800 42498 10540 42530
rect 9800 1000 10100 42498
rect 14130 42470 14550 42480
rect 14130 42370 14140 42470
rect 14240 42468 14550 42470
rect 14240 42370 27016 42468
rect 14130 42360 27016 42370
rect 14548 42348 27016 42360
rect 400 0 520 200
rect 4816 0 4936 200
rect 9232 0 9352 200
rect 13648 0 13768 200
rect 18064 0 18184 200
rect 22480 0 22600 200
rect 26896 0 27016 42348
rect 31318 34278 31426 43004
rect 31319 200 31425 34278
rect 31312 0 31432 200
<< labels >>
flabel metal4 s 30974 44952 31034 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 31710 44952 31770 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 30238 44952 30298 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 31312 0 31432 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26896 0 27016 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22480 0 22600 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18064 0 18184 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 13648 0 13768 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 9232 0 9352 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 4816 0 4936 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 400 0 520 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 29502 44952 29562 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 28030 44952 28090 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 27294 44952 27354 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 25822 44952 25882 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 25086 44952 25146 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23614 44952 23674 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22878 44952 22938 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21406 44952 21466 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 20670 44952 20730 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19198 44952 19258 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 18462 44952 18522 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 5950 44952 6010 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 5214 44952 5274 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 4478 44952 4538 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 3742 44952 3802 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 3006 44952 3066 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 2270 44952 2330 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 1534 44952 1594 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 798 44952 858 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 10366 44952 10426 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 9630 44952 9690 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 8158 44952 8218 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 7422 44952 7482 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 16990 44952 17050 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 16254 44952 16314 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 14782 44952 14842 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 14046 44952 14106 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 12574 44952 12634 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 11838 44952 11898 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 200 1000 500 44152 1 FreeSans 2 0 0 0 VPWR
port 51 nsew power bidirectional
rlabel locali 13510 42880 13550 42920 1 Y
rlabel locali 13250 42920 13290 42960 1 A
flabel metal4 9800 1000 10100 44152 1 FreeSans 2 0 0 0 VGND
port 52 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
