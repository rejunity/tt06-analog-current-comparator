* NGSPICE file created from tt_um_rejunity_current_cmp.ext - technology: sky130A

 clk ena rst_n ua[0] ua[1] ua[2] ua[3] ua[4] ua[5]
+ ua[6] ua[7] ui_in[0] ui_in[1] ui_in[2] ui_in[3] ui_in[4] ui_in[5] ui_in[6] ui_in[7]
+ uio_in[0] uio_in[1] uio_in[2] uio_in[3] uio_in[4] uio_in[5] uio_in[6] uio_in[7]
+ VPWR VGND
X0 a_21880_41750# a_21880_41750# VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.35 pd=2.7 as=0.4 ps=2.8 w=1 l=0.15
X1 a_21880_41750# a_22050_41640# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.54 as=0.168 ps=1.64 w=0.42 l=0.15
R0 uio_in[0] a_23490_41640# sky130_fd_pr__res_generic_m2 w=0.45 l=0.05
X2 a_21880_41750# a_22530_41640# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.54 as=0.168 ps=1.64 w=0.42 l=0.15
X3 a_24200_41490# a_24200_41490# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.54 as=0.168 ps=1.64 w=0.42 l=0.15
X4 a_24200_41490# a_25370_41750# VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.35 pd=2.7 as=0.4 ps=2.8 w=1 l=0.15
X5 a_23810_40680# Idiff VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.45 pd=2.9 as=0.4 ps=2.8 w=1 l=0.15
X6 a_24200_41490# a_25850_41750# VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.35 pd=2.7 as=0.4 ps=2.8 w=1 l=0.15
X7 a_24200_41490# a_24410_41750# VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.35 pd=2.7 as=0.4 ps=2.8 w=1 l=0.15
X8 a_24200_41490# a_24200_41490# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.54 as=0.168 ps=1.64 w=0.42 l=0.15
X9 a_23810_40680# Idiff VGND VGND sky130_fd_pr__nfet_01v8 ad=0.189 pd=1.74 as=0.168 ps=1.64 w=0.42 l=0.15
X10 a_13070_38680# a_13100_38710# w_12870_38970# w_12870_38970# sky130_fd_pr__pfet_01v8 ad=0.45 pd=2.9 as=0.4 ps=2.8 w=1 l=0.15
X11 a_24200_41490# a_24890_41750# VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.35 pd=2.7 as=0.4 ps=2.8 w=1 l=0.15
X12 a_24200_41490# a_24200_41490# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.54 as=0.168 ps=1.64 w=0.42 l=0.15
X13 a_24200_41490# a_24200_41490# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.54 as=0.168 ps=1.64 w=0.42 l=0.15
R1 uio_in[5] a_22290_41640# sky130_fd_pr__res_generic_m2 w=0.45 l=0.05
X14 a_24200_41490# a_24200_41490# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.54 as=0.168 ps=1.64 w=0.42 l=0.15
X15 Idiff a_23810_40680# VGND VPWR sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.8 ps=3.6 w=1 l=0.15
X16 a_13070_38680# a_13100_38710# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.189 pd=1.74 as=0.168 ps=1.64 w=0.42 l=0.15
X17 a_24200_41490# a_25130_41750# VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.35 pd=2.7 as=0.4 ps=2.8 w=1 l=0.15
X18 Idiff a_23810_40680# VPWR VGND sky130_fd_pr__nfet_01v8 ad=0.168 pd=1.64 as=0.189 ps=1.74 w=0.42 l=0.15
X19 VGND a_24200_41490# Idiff VGND sky130_fd_pr__nfet_01v8 ad=0.231 pd=1.94 as=0.231 ps=1.94 w=0.42 l=0.15
X20 a_24200_41490# a_24200_41490# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.54 as=0.168 ps=1.64 w=0.42 l=0.15
X21 a_24200_41490# a_24650_41750# VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.35 pd=2.7 as=0.4 ps=2.8 w=1 l=0.15
X22 a_24200_41490# a_24200_41490# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.54 as=0.168 ps=1.64 w=0.42 l=0.15
R2 uio_in[2] a_23010_41640# sky130_fd_pr__res_generic_m2 w=0.45 l=0.05
R3 ui_in[2] a_25610_41750# sky130_fd_pr__res_generic_m2 w=0.45 l=0.05
R4 ui_in[6] a_24650_41750# sky130_fd_pr__res_generic_m2 w=0.45 l=0.05
X23 a_21880_41750# a_21880_41750# VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.35 pd=2.7 as=0.4 ps=2.8 w=1 l=0.15
X24 a_21880_41750# a_21880_41750# VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.35 pd=2.7 as=0.4 ps=2.8 w=1 l=0.15
R5 ui_in[3] a_25370_41750# sky130_fd_pr__res_generic_m2 w=0.45 l=0.05
X25 a_21880_41750# a_23010_41640# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.54 as=0.168 ps=1.64 w=0.42 l=0.15
R6 ui_in[7] a_24410_41750# sky130_fd_pr__res_generic_m2 w=0.45 l=0.05
X26 a_21880_41750# a_23490_41640# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.54 as=0.168 ps=1.64 w=0.42 l=0.15
R7 uio_in[3] a_22770_41640# sky130_fd_pr__res_generic_m2 w=0.45 l=0.05
R8 uio_in[4] a_22530_41640# sky130_fd_pr__res_generic_m2 w=0.45 l=0.05
X27 a_21880_41750# a_21880_41750# VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.35 pd=2.7 as=0.4 ps=2.8 w=1 l=0.15
X28 a_21880_41750# a_23250_41640# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.54 as=0.168 ps=1.64 w=0.42 l=0.15
R9 ui_in[4] a_25130_41750# sky130_fd_pr__res_generic_m2 w=0.45 l=0.05
R10 ui_in[0] a_26090_41750# sky130_fd_pr__res_generic_m2 w=0.45 l=0.05
X29 a_21880_41750# a_21880_41750# VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.35 pd=2.7 as=0.4 ps=2.8 w=1 l=0.15
X30 ua[0] a_23810_40680# VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.45 pd=2.9 as=0.4 ps=2.8 w=1 l=0.15
X31 a_21880_41750# a_21880_41750# VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.35 pd=2.7 as=0.4 ps=2.8 w=1 l=0.15
X32 Idiff a_21880_41750# VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.55 pd=3.1 as=0.55 ps=3.1 w=1 l=0.15
X33 a_21880_41750# a_22290_41640# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.54 as=0.168 ps=1.64 w=0.42 l=0.15
X34 a_13100_38710# a_13070_38680# VGND w_12870_38970# sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.8 ps=3.6 w=1 l=0.15
X35 a_21880_41750# a_21880_41750# VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.35 pd=2.7 as=0.4 ps=2.8 w=1 l=0.15
X36 a_21880_41750# a_22770_41640# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.54 as=0.168 ps=1.64 w=0.42 l=0.15
R11 uio_in[6] a_22050_41640# sky130_fd_pr__res_generic_m2 w=0.45 l=0.05
R12 ui_in[5] a_24890_41750# sky130_fd_pr__res_generic_m2 w=0.45 l=0.05
X37 a_24200_41490# a_26090_41750# VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.35 pd=2.7 as=0.4 ps=2.8 w=1 l=0.15
X38 ua[0] a_23810_40680# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.189 pd=1.74 as=0.168 ps=1.64 w=0.42 l=0.15
X39 a_13100_38710# a_13070_38680# w_12870_38970# VGND sky130_fd_pr__nfet_01v8 ad=0.168 pd=1.64 as=0.189 ps=1.74 w=0.42 l=0.15
R13 uio_in[1] a_23250_41640# sky130_fd_pr__res_generic_m2 w=0.45 l=0.05
X40 a_21880_41750# a_21810_41640# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.54 as=0.168 ps=1.64 w=0.42 l=0.15
X41 a_24200_41490# a_24200_41490# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.54 as=0.168 ps=1.64 w=0.42 l=0.15
X42 a_21880_41750# a_21880_41750# VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.35 pd=2.7 as=0.4 ps=2.8 w=1 l=0.15
X43 a_24200_41490# a_25610_41750# VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.35 pd=2.7 as=0.4 ps=2.8 w=1 l=0.15
R14 uio_in[7] a_21810_41640# sky130_fd_pr__res_generic_m2 w=0.45 l=0.05
R15 ui_in[1] a_25850_41750# sky130_fd_pr__res_generic_m2 w=0.45 l=0.05
C0 m2_21390_44110# m2_22130_44110# 0.007143f
C1 m2_20650_44110# m2_21390_44110# 0.007143f
C2 m2_19910_44110# m2_20650_44110# 0.007143f
C3 clk ena 0.023797f
C4 w_12870_38970# m1_13270_38360# 0.00635f
C5 m2_19170_44110# m2_19910_44110# 0.007143f
C6 rst_n clk 0.023797f
C7 m2_18430_44110# m2_19170_44110# 0.007143f
C8 ui_in[0] rst_n 0.023797f
C9 ui_in[1] ui_in[0] 0.13387f
C10 ui_in[2] ui_in[1] 0.133768f
C11 ui_in[3] ui_in[2] 0.133458f
C12 ui_in[4] ui_in[3] 0.133435f
C13 ui_in[5] ui_in[4] 0.133252f
C14 ui_in[6] ui_in[5] 0.133228f
C15 ui_in[7] ui_in[6] 0.13321f
C16 VPWR ua[7] 0.010285f
C17 uio_in[0] ui_in[7] 0.132332f
C18 a_13100_38710# li_14140_38880# 0.008859f
C19 a_13070_38680# li_14140_38880# 0.011142f
C20 uio_in[1] uio_in[0] 0.134137f
C21 a_13070_38680# a_13100_38710# 0.250071f
C22 uio_in[2] uio_in[1] 0.13321f
C23 a_23490_41640# uio_in[0] 0.044617f
C24 m2_29530_44110# ui_in[0] 0.020029f
C25 uio_in[3] uio_in[2] 0.13321f
C26 a_23250_41640# uio_in[1] 0.043751f
C27 a_26090_41750# ui_in[0] 0.049656f
C28 VPWR ui_in[4] 0.004568f
C29 m2_28790_44110# ui_in[1] 0.020255f
C30 a_26090_41750# ui_in[1] 3.52e-19
C31 a_23010_41640# uio_in[1] 0.001582f
C32 VPWR ui_in[5] 0.004568f
C33 uio_in[4] uio_in[3] 0.13321f
C34 a_25850_41750# ui_in[1] 0.049419f
C35 a_26090_41750# ui_in[2] 3.3e-19
C36 a_23010_41640# uio_in[2] 0.046102f
C37 a_23250_41640# a_23490_41640# 0.473575f
C38 VPWR ui_in[6] 0.004568f
C39 m2_28050_44110# ui_in[2] 0.02048f
C40 a_25850_41750# ui_in[2] 5.76e-19
C41 a_26090_41750# ui_in[3] 3.3e-19
C42 a_22770_41640# uio_in[2] 0.001135f
C43 VPWR ui_in[7] 0.004568f
C44 uio_in[5] uio_in[4] 0.13321f
C45 a_25610_41750# ui_in[2] 0.051252f
C46 a_25850_41750# ui_in[3] 5.66e-19
C47 a_26090_41750# ui_in[4] 3.3e-19
C48 a_22530_41640# uio_in[2] 8.23e-19
C49 a_22770_41640# uio_in[3] 0.047856f
C50 a_23010_41640# a_23250_41640# 0.526351f
C51 VPWR uio_in[0] 0.004568f
C52 m2_27310_44110# ui_in[3] 0.020706f
C53 a_25610_41750# ui_in[3] 6.72e-19
C54 a_25850_41750# ui_in[4] 5.53e-19
C55 a_22290_41640# uio_in[2] 6.38e-19
C56 a_22530_41640# uio_in[3] 8.23e-19
C57 VPWR uio_in[1] 0.004568f
C58 uio_in[6] uio_in[5] 0.13321f
C59 a_22530_41640# uio_in[4] 0.049358f
C60 a_25370_41750# ui_in[3] 0.049254f
C61 a_25610_41750# ui_in[4] 6.57e-19
C62 a_23810_40680# ua[0] 0.067902f
C63 a_25850_41750# ui_in[5] 0.001163f
C64 a_22290_41640# uio_in[3] 6.38e-19
C65 a_22770_41640# a_23010_41640# 0.642783f
C66 VPWR uio_in[2] 0.004568f
C67 m2_26570_44110# ui_in[4] 0.020932f
C68 a_22050_41640# uio_in[3] 5.15e-19
C69 a_22290_41640# uio_in[4] 6.38e-19
C70 a_25370_41750# ui_in[4] 8.82e-19
C71 a_25610_41750# ui_in[5] 6.45e-19
C72 a_23810_40680# VPWR 0.250758f
C73 a_22530_41640# a_23010_41640# 1.6e-19
C74 VPWR uio_in[3] 0.004568f
C75 uio_in[7] uio_in[6] 0.13321f
C76 a_22050_41640# uio_in[4] 5.15e-19
C77 a_22290_41640# uio_in[5] 0.050403f
C78 a_25370_41750# ui_in[5] 8.67e-19
C79 a_21810_41640# uio_in[3] 2.96e-19
C80 a_23490_41640# VPWR 0.272141f
C81 a_25130_41750# ui_in[4] 0.048012f
C82 a_22290_41640# a_23010_41640# 1.13e-19
C83 a_22530_41640# a_22770_41640# 0.720865f
C84 a_24200_41490# a_23810_40680# 0.001209f
C85 m2_25830_44110# ui_in[5] 0.021157f
C86 VPWR uio_in[4] 0.004568f
C87 a_22050_41640# uio_in[5] 5.15e-19
C88 a_21810_41640# uio_in[4] 2.96e-19
C89 a_23250_41640# VPWR 0.225848f
C90 a_25130_41750# ui_in[5] 0.001175f
C91 a_22290_41640# a_22770_41640# 1.23e-19
C92 Idiff a_23810_40680# 0.274331f
C93 a_24200_41490# a_23490_41640# 0.004679f
C94 a_22050_41640# uio_in[6] 0.051224f
C95 a_21810_41640# uio_in[5] 2.96e-19
C96 a_23010_41640# VPWR 0.22923f
C97 a_24890_41750# ui_in[5] 0.046777f
C98 a_25130_41750# ui_in[6] 0.004014f
C99 a_22290_41640# a_22530_41640# 0.900719f
C100 a_22050_41640# a_22770_41640# 9.52e-20
C101 a_24200_41490# a_23250_41640# 1.08e-20
C102 Idiff a_23490_41640# 0.005611f
C103 m2_25090_44110# ui_in[6] 0.021383f
C104 a_24890_41750# ui_in[6] 0.001608f
C105 a_21810_41640# uio_in[6] 2.96e-19
C106 a_22770_41640# VPWR 0.235182f
C107 a_22050_41640# a_22530_41640# 1.18e-19
C108 Idiff a_23250_41640# 2.72e-19
C109 a_24200_41490# a_23010_41640# 6.92e-21
C110 a_21810_41640# a_22770_41640# 7.47e-20
C111 a_24650_41750# ui_in[6] 0.044593f
C112 a_21810_41640# uio_in[7] 0.050442f
C113 a_22530_41640# VPWR 0.248503f
C114 a_22050_41640# a_22290_41640# 1.08768f
C115 Idiff a_23010_41640# 1.47e-19
C116 a_24200_41490# a_22770_41640# 4.79e-21
C117 a_21810_41640# a_22530_41640# 9.71e-20
C118 m2_24350_44110# ui_in[7] 0.021608f
C119 a_22290_41640# VPWR 0.266254f
C120 Idiff a_22770_41640# 9.1e-20
C121 a_24200_41490# a_22530_41640# 4.57e-22
C122 a_21810_41640# a_22290_41640# 1.06e-19
C123 VPWR ua[0] 0.499805f
C124 a_24410_41750# ui_in[7] 0.044373f
C125 a_22050_41640# VPWR 0.297591f
C126 Idiff a_22530_41640# 6.16e-20
C127 a_21810_41640# a_22050_41640# 1.10845f
C128 m2_23590_44110# uio_in[0] 0.021608f
C129 a_21810_41640# VPWR 0.61255f
C130 a_24200_41490# ua[0] 0.020222f
C131 Idiff a_22290_41640# 4.44e-20
C132 a_24200_41490# VPWR 1.32326f
C133 Idiff ua[0] 0.007155f
C134 w_12870_38970# li_14140_38880# 0.00761f
C135 m2_22870_44110# uio_in[1] 0.021608f
C136 Idiff VPWR 0.591003f
C137 a_26090_41750# ua[0] 0.003257f
C138 w_12870_38970# a_13100_38710# 0.411194f
C139 a_24410_41750# a_23810_40680# 0.001267f
C140 a_26090_41750# VPWR 0.510899f
C141 a_25850_41750# ua[0] 0.003181f
C142 a_23490_41640# m2_23590_44110# 0.005112f
C143 Idiff a_24200_41490# 0.02177f
C144 w_12870_38970# a_13070_38680# 0.147772f
C145 a_24410_41750# a_23490_41640# 0.128679f
C146 a_21880_41750# a_23810_40680# 0.002387f
C147 m2_22130_44110# uio_in[2] 0.021608f
C148 a_25850_41750# VPWR 0.317633f
C149 a_25610_41750# ua[0] 0.003257f
C150 a_26090_41750# a_24200_41490# 0.14468f
C151 a_21880_41750# a_23490_41640# 0.212873f
C152 m2_28790_44110# m2_29530_44110# 0.007143f
C153 a_25610_41750# VPWR 0.306437f
C154 a_25370_41750# ua[0] 0.003295f
C155 a_23250_41640# m2_22870_44110# 0.005112f
C156 a_26090_41750# m2_29530_44110# 0.005112f
C157 a_25850_41750# a_24200_41490# 0.144319f
C158 a_21880_41750# a_23250_41640# 0.204944f
C159 m2_21390_44110# uio_in[3] 0.021608f
C160 a_25370_41750# VPWR 0.29637f
C161 a_25130_41750# ua[0] 0.002253f
C162 a_25610_41750# a_24200_41490# 0.144119f
C163 a_21880_41750# a_23010_41640# 0.205094f
C164 m2_28050_44110# m2_28790_44110# 0.007143f
C165 a_25850_41750# m2_28790_44110# 0.005112f
C166 a_24890_41750# ua[0] 8.21e-20
C167 a_23010_41640# m2_22130_44110# 0.005112f
C168 li_14140_38880# m1_13270_38360# 0.057421f
C169 a_25130_41750# VPWR 0.288147f
C170 a_25370_41750# a_24200_41490# 0.143902f
C171 a_25850_41750# a_26090_41750# 1.12631f
C172 a_21880_41750# a_22770_41640# 0.205425f
C173 m2_20650_44110# uio_in[4] 0.021608f
C174 a_13100_38710# m1_13270_38360# 0.0037f
C175 a_24890_41750# VPWR 0.278208f
C176 a_24650_41750# ua[0] 1.32e-19
C177 a_25130_41750# a_24200_41490# 0.143584f
C178 a_25610_41750# a_26090_41750# 1.54e-19
C179 a_21880_41750# a_22530_41640# 0.205638f
C180 m2_27310_44110# m2_28050_44110# 0.007143f
C181 a_13070_38680# m1_13270_38360# 0.005568f
C182 a_24650_41750# VPWR 0.265643f
C183 a_25610_41750# m2_28050_44110# 0.005112f
C184 a_24410_41750# ua[0] 0.001226f
C185 a_22770_41640# m2_21390_44110# 0.005112f
C186 a_24890_41750# a_24200_41490# 0.143416f
C187 a_25370_41750# a_26090_41750# 1.28e-19
C188 a_25610_41750# a_25850_41750# 1.33939f
C189 a_21880_41750# a_22290_41640# 0.205822f
C190 m2_19910_44110# uio_in[5] 0.021608f
C191 a_24410_41750# VPWR 0.316454f
C192 a_24650_41750# a_24200_41490# 0.1433f
C193 a_25130_41750# a_26090_41750# 1.13e-19
C194 a_25370_41750# a_25850_41750# 1.49e-19
C195 a_21880_41750# a_22050_41640# 0.206073f
C196 m2_26570_44110# m2_27310_44110# 0.007143f
C197 a_22530_41640# m2_20650_44110# 0.005112f
C198 a_21880_41750# VPWR 1.67321f
C199 a_25370_41750# m2_27310_44110# 0.005112f
C200 a_24410_41750# a_24200_41490# 0.111243f
C201 a_25130_41750# a_25850_41750# 1.34e-19
C202 a_21880_41750# a_21810_41640# 0.159038f
C203 a_25370_41750# a_25610_41750# 0.812521f
C204 m2_19170_44110# uio_in[6] 0.021608f
C205 a_21880_41750# a_24200_41490# 0.001258f
C206 a_24410_41750# Idiff 0.007045f
C207 a_24890_41750# a_25850_41750# 3.05e-19
C208 a_25130_41750# a_25610_41750# 1.56e-19
C209 m2_25830_44110# m2_26570_44110# 0.007143f
C210 a_22290_41640# m2_19910_44110# 0.005112f
C211 a_25130_41750# m2_26570_44110# 0.005112f
C212 a_21880_41750# Idiff 0.072467f
C213 a_24890_41750# a_25610_41750# 1.23e-19
C214 a_25130_41750# a_25370_41750# 0.758603f
C215 m2_18430_44110# uio_in[7] 0.021608f
C216 a_24890_41750# a_25370_41750# 1.78e-19
C217 m2_25090_44110# m2_25830_44110# 0.007143f
C218 a_22050_41640# m2_19170_44110# 0.005112f
C219 a_24890_41750# m2_25830_44110# 0.005112f
C220 a_24890_41750# a_25130_41750# 0.652808f
C221 a_24650_41750# a_25130_41750# 8.46e-19
C222 m2_24350_44110# m2_25090_44110# 0.007143f
C223 a_24650_41750# m2_25090_44110# 0.005112f
C224 a_21810_41640# m2_18430_44110# 0.005112f
C225 a_21880_41750# a_25370_41750# 4.13e-21
C226 a_24650_41750# a_24890_41750# 0.550955f
C227 a_21880_41750# a_25130_41750# 5.8e-21
C228 m2_23590_44110# m2_24350_44110# 0.006944f
C229 a_24410_41750# m2_24350_44110# 0.005112f
C230 a_21880_41750# a_24890_41750# 8.71e-21
C231 a_24410_41750# a_24650_41750# 0.454394f
C232 a_21880_41750# a_24650_41750# 1.44e-20
C233 m2_22870_44110# m2_23590_44110# 0.007353f
C234 a_21880_41750# a_24410_41750# 0.006714f
C235 m2_22130_44110# m2_22870_44110# 0.007143f
C236 ua[2] VGND 0.122428f
C237 ua[3] VGND 0.122428f
C238 ua[4] VGND 0.122428f
C239 ua[5] VGND 0.122428f
C240 ua[6] VGND 0.122428f
C241 ua[7] VGND 0.111009f
C242 ena VGND 0.073297f
C243 clk VGND 0.0487f
C244 rst_n VGND 0.0487f
C245 ui_in[0] VGND 0.350951f
C246 ui_in[1] VGND 0.234234f
C247 ui_in[2] VGND 0.230502f
C248 ui_in[3] VGND 0.230704f
C249 ui_in[4] VGND 0.223397f
C250 ui_in[5] VGND 0.22191f
C251 ui_in[6] VGND 0.220814f
C252 ui_in[7] VGND 0.223871f
C253 uio_in[0] VGND 0.225466f
C254 uio_in[1] VGND 0.224179f
C255 uio_in[2] VGND 0.221286f
C256 uio_in[3] VGND 0.219592f
C257 uio_in[4] VGND 0.218871f
C258 uio_in[5] VGND 0.224716f
C259 uio_in[6] VGND 0.224366f
C260 uio_in[7] VGND 0.362103f
C261 ua[1] VGND 16.757198f
C262 ua[0] VGND 18.8739f
C263 VPWR VGND 53.1585f
C264 m2_29530_44110# VGND 0.049454f $ **FLOATING
C265 m2_28790_44110# VGND 0.040694f $ **FLOATING
C266 m2_28050_44110# VGND 0.040694f $ **FLOATING
C267 m2_27310_44110# VGND 0.040694f $ **FLOATING
C268 m2_26570_44110# VGND 0.040694f $ **FLOATING
C269 m2_25830_44110# VGND 0.040694f $ **FLOATING
C270 m2_25090_44110# VGND 0.040694f $ **FLOATING
C271 m2_24350_44110# VGND 0.040877f $ **FLOATING
C272 m2_23590_44110# VGND 0.040687f $ **FLOATING
C273 m2_22870_44110# VGND 0.040504f $ **FLOATING
C274 m2_22130_44110# VGND 0.040694f $ **FLOATING
C275 m2_21390_44110# VGND 0.040694f $ **FLOATING
C276 m2_20650_44110# VGND 0.040694f $ **FLOATING
C277 m2_19910_44110# VGND 0.040694f $ **FLOATING
C278 m2_19170_44110# VGND 0.040694f $ **FLOATING
C279 m2_18430_44110# VGND 0.049454f $ **FLOATING
C280 m1_13270_38360# VGND 0.934988f $ **FLOATING
C281 li_14140_38880# VGND 0.665446f $ **FLOATING
C282 a_13100_38710# VGND 0.453185f
C283 a_13070_38680# VGND 0.542482f
C284 a_23810_40680# VGND 0.717709f
C285 a_23490_41640# VGND 0.839973f
C286 a_23250_41640# VGND 0.763056f
C287 a_23010_41640# VGND 0.903577f
C288 a_22770_41640# VGND 1.00469f
C289 a_22530_41640# VGND 1.09077f
C290 a_22290_41640# VGND 1.16005f
C291 a_22050_41640# VGND 1.25686f
C292 a_21810_41640# VGND 2.12497f
C293 a_24200_41490# VGND 2.65987f
C294 Idiff VGND 0.750117f
C295 a_26090_41750# VGND 1.99112f
C296 a_25850_41750# VGND 1.14437f
C297 a_25610_41750# VGND 1.06238f
C298 a_25370_41750# VGND 1.02102f
C299 a_25130_41750# VGND 0.909708f
C300 a_24890_41750# VGND 0.808573f
C301 a_24650_41750# VGND 0.69159f
C302 a_24410_41750# VGND 0.702523f
C303 a_21880_41750# VGND 1.94325f
C304 w_12870_38970# VGND 1.34935f


