.ends

* set gnd and power
Vgnd VGND 0 0
Vdd VPWR VGND 1.8

* create pulse
* Vin A VGND pulse(0 1.8 1p 10p 10p 1n 2n)
* Isource A VGND pulse(-0.001 0.001 0 500p 500p 500p 2n)

* Vin0 X0 VGND pulse(0 1.8 1p 10p 10p 1n 2n)
* Vin1 X1 VGND 0
* Vin2 Y0 VGND pulse(0 1.8 500p 10p 10p 1n 2n)
* Vin3 Y1 VGND 0
* .tran 10e-12 2e-09 0e-00

*   112233
*  5050505
* 01210121
* 000011112222

* pulse(0 1.8  5n 10p 10p 10n 20n)
* pulse(0 1.8 10n 10p 10p 10n 20n)
* pulse(0 1.8 20n 10p 10p 20n 40n)
* pulse(0 1.8  1p 10p 10p 20n 40n)

Vin0 X0 VGND pulse(1.8 0 20n 10p 10p 40n 80n)
Vin1 X1 VGND pulse(1.8 0 40n 10p 10p 40n 80n)
Vin2 Y0 VGND pulse(0 1.8  5n 10p 10p 10n 20n)
Vin3 Y1 VGND pulse(0 1.8 10n 10p 10p 10n 20n)
.tran 10e-12 6e-08 0e-00

.control
run
set color0 = white
set color1 = black
plot X0, X1
plot Y0, Y1
plot Out
plot i(Vdd)
.endc