* NGSPICE file created from tt_um_rejunity_current_cmp.ext - technology: sky130A

 clk ena rst_n ua[0] ua[2] ua[3] ua[4] ua[5] ua[6]
+ ua[7] ui_in[0] ui_in[1] ui_in[2] ui_in[3] ui_in[4] ui_in[5] ui_in[6] ui_in[7] uio_in[0]
+ uio_in[1] uio_in[2] uio_in[3] uio_in[4] uio_in[5] uio_in[6] uio_in[7] VPWR VGND
+ ua[1]
X0 a_21880_41750# a_21880_41750# VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.35 pd=2.7 as=0.4 ps=2.8 w=1 l=0.15
X1 a_21880_41750# a_22050_39050# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.54 as=0.168 ps=1.64 w=0.42 l=0.15
R0 uio_in[0] a_23490_39050# sky130_fd_pr__res_generic_m2 w=0.45 l=0.05
X2 a_21880_41750# a_22530_39050# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.54 as=0.168 ps=1.64 w=0.42 l=0.15
X3 a_24200_41490# a_24200_41490# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.54 as=0.168 ps=1.64 w=0.42 l=0.15
X4 a_21880_39160# a_21880_39160# VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.35 pd=2.7 as=0.4 ps=2.8 w=1 l=0.15
X5 a_21880_39160# a_22050_39050# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.54 as=0.168 ps=1.64 w=0.42 l=0.15
X6 a_21880_39160# a_21880_39160# VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.35 pd=2.7 as=0.4 ps=2.8 w=1 l=0.15
X7 a_24200_38900# a_25610_39160# VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.35 pd=2.7 as=0.4 ps=2.8 w=1 l=0.15
X8 a_21880_39160# a_22530_39050# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.54 as=0.168 ps=1.64 w=0.42 l=0.15
X9 a_24200_38900# a_24200_38900# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.54 as=0.168 ps=1.64 w=0.42 l=0.15
X10 a_24200_41490# a_25370_39160# VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.35 pd=2.7 as=0.4 ps=2.8 w=1 l=0.15
X11 a_23810_40680# ua[1] VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.45 pd=2.9 as=0.4 ps=2.8 w=1 l=0.15
X12 a_24200_41490# a_25850_39160# VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.35 pd=2.7 as=0.4 ps=2.8 w=1 l=0.15
X13 a_24200_41490# a_24410_39160# VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.35 pd=2.7 as=0.4 ps=2.8 w=1 l=0.15
X14 a_24200_41490# a_24200_41490# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.54 as=0.168 ps=1.64 w=0.42 l=0.15
X15 a_23810_40680# ua[1] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.189 pd=1.74 as=0.168 ps=1.64 w=0.42 l=0.15
X16 a_13070_38680# a_13100_38710# w_12870_38970# w_12870_38970# sky130_fd_pr__pfet_01v8 ad=0.45 pd=2.9 as=0.4 ps=2.8 w=1 l=0.15
X17 a_24200_41490# a_24890_39160# VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.35 pd=2.7 as=0.4 ps=2.8 w=1 l=0.15
X18 a_24200_41490# a_24200_41490# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.54 as=0.168 ps=1.64 w=0.42 l=0.15
X19 a_24200_41490# a_24200_41490# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.54 as=0.168 ps=1.64 w=0.42 l=0.15
X20 a_24200_38900# a_25370_39160# VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.35 pd=2.7 as=0.4 ps=2.8 w=1 l=0.15
X21 a_24200_38900# a_24200_38900# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.54 as=0.168 ps=1.64 w=0.42 l=0.15
R1 uio_in[5] a_22290_39050# sky130_fd_pr__res_generic_m2 w=0.45 l=0.05
X22 a_24200_41490# a_24200_41490# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.54 as=0.168 ps=1.64 w=0.42 l=0.15
X23 ua[1] a_23810_40680# VGND VPWR sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.8 ps=3.6 w=1 l=0.15
X24 a_24200_38900# a_25850_39160# VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.35 pd=2.7 as=0.4 ps=2.8 w=1 l=0.15
X25 a_24200_38900# a_24200_38900# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.54 as=0.168 ps=1.64 w=0.42 l=0.15
X26 a_24200_38900# a_24200_38900# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.54 as=0.168 ps=1.64 w=0.42 l=0.15
X27 a_13070_38680# a_13100_38710# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.189 pd=1.74 as=0.168 ps=1.64 w=0.42 l=0.15
X28 a_24200_41490# a_25130_39160# VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.35 pd=2.7 as=0.4 ps=2.8 w=1 l=0.15
X29 a_24200_38900# a_24410_39160# VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.35 pd=2.7 as=0.4 ps=2.8 w=1 l=0.15
X30 a_24200_38900# a_24200_38900# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.54 as=0.168 ps=1.64 w=0.42 l=0.15
X31 ua[1] a_23810_40680# VPWR VGND sky130_fd_pr__nfet_01v8 ad=0.168 pd=1.64 as=0.189 ps=1.74 w=0.42 l=0.15
X32 a_24200_38900# a_24890_39160# VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.35 pd=2.7 as=0.4 ps=2.8 w=1 l=0.15
X33 VGND a_24200_41490# ua[1] VGND sky130_fd_pr__nfet_01v8 ad=0.231 pd=1.94 as=0.231 ps=1.94 w=0.42 l=0.15
X34 a_24200_41490# a_24200_41490# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.54 as=0.168 ps=1.64 w=0.42 l=0.15
X35 a_24200_41490# a_24650_39160# VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.35 pd=2.7 as=0.4 ps=2.8 w=1 l=0.15
X36 a_24200_38900# a_25130_39160# VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.35 pd=2.7 as=0.4 ps=2.8 w=1 l=0.15
X37 VGND a_24200_38900# ua[1] VGND sky130_fd_pr__nfet_01v8 ad=0.231 pd=1.94 as=0.231 ps=1.94 w=0.42 l=0.15
X38 a_24200_38900# a_24200_38900# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.54 as=0.168 ps=1.64 w=0.42 l=0.15
X39 a_24200_41490# a_24200_41490# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.54 as=0.168 ps=1.64 w=0.42 l=0.15
X40 a_24200_38900# a_24650_39160# VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.35 pd=2.7 as=0.4 ps=2.8 w=1 l=0.15
X41 a_24200_38900# a_24200_38900# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.54 as=0.168 ps=1.64 w=0.42 l=0.15
R2 uio_in[2] a_23010_39050# sky130_fd_pr__res_generic_m2 w=0.45 l=0.05
R3 ui_in[2] a_25610_39160# sky130_fd_pr__res_generic_m2 w=0.45 l=0.05
R4 ui_in[6] a_24650_39160# sky130_fd_pr__res_generic_m2 w=0.45 l=0.05
X42 a_21880_41750# a_21880_41750# VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.35 pd=2.7 as=0.4 ps=2.8 w=1 l=0.15
X43 a_21880_41750# a_21880_41750# VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.35 pd=2.7 as=0.4 ps=2.8 w=1 l=0.15
R5 ui_in[3] a_25370_39160# sky130_fd_pr__res_generic_m2 w=0.45 l=0.05
X44 a_21880_41750# a_23010_39050# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.54 as=0.168 ps=1.64 w=0.42 l=0.15
R6 ui_in[7] a_24410_39160# sky130_fd_pr__res_generic_m2 w=0.45 l=0.05
X45 a_21880_41750# a_23490_39050# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.54 as=0.168 ps=1.64 w=0.42 l=0.15
X46 a_21880_39160# a_21880_39160# VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.35 pd=2.7 as=0.4 ps=2.8 w=1 l=0.15
X47 a_21880_39160# a_23010_39050# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.54 as=0.168 ps=1.64 w=0.42 l=0.15
R7 uio_in[3] a_22770_39050# sky130_fd_pr__res_generic_m2 w=0.45 l=0.05
X48 a_21880_39160# a_21880_39160# VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.35 pd=2.7 as=0.4 ps=2.8 w=1 l=0.15
X49 a_21880_39160# a_23490_39050# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.54 as=0.168 ps=1.64 w=0.42 l=0.15
R8 uio_in[4] a_22530_39050# sky130_fd_pr__res_generic_m2 w=0.45 l=0.05
X50 a_21880_41750# a_21880_41750# VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.35 pd=2.7 as=0.4 ps=2.8 w=1 l=0.15
X51 a_21880_41750# a_23250_39050# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.54 as=0.168 ps=1.64 w=0.42 l=0.15
R9 ui_in[4] a_25130_39160# sky130_fd_pr__res_generic_m2 w=0.45 l=0.05
R10 ui_in[0] a_26090_39160# sky130_fd_pr__res_generic_m2 w=0.45 l=0.05
X52 a_21880_41750# a_21880_41750# VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.35 pd=2.7 as=0.4 ps=2.8 w=1 l=0.15
X53 ua[0] a_23810_40680# VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.45 pd=2.9 as=0.4 ps=2.8 w=1 l=0.15
X54 a_21880_41750# a_21880_41750# VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.35 pd=2.7 as=0.4 ps=2.8 w=1 l=0.15
X55 ua[1] a_21880_41750# VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.55 pd=3.1 as=0.55 ps=3.1 w=1 l=0.15
X56 a_21880_41750# a_22290_39050# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.54 as=0.168 ps=1.64 w=0.42 l=0.15
X57 a_21880_39160# a_21880_39160# VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.35 pd=2.7 as=0.4 ps=2.8 w=1 l=0.15
X58 a_13100_38710# a_13070_38680# VGND w_12870_38970# sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.8 ps=3.6 w=1 l=0.15
X59 a_21880_39160# a_23250_39050# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.54 as=0.168 ps=1.64 w=0.42 l=0.15
X60 a_21880_41750# a_21880_41750# VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.35 pd=2.7 as=0.4 ps=2.8 w=1 l=0.15
X61 a_21880_41750# a_22770_39050# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.54 as=0.168 ps=1.64 w=0.42 l=0.15
X62 a_21880_39160# a_21880_39160# VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.35 pd=2.7 as=0.4 ps=2.8 w=1 l=0.15
X63 a_21880_39160# a_22290_39050# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.54 as=0.168 ps=1.64 w=0.42 l=0.15
R11 uio_in[6] a_22050_39050# sky130_fd_pr__res_generic_m2 w=0.45 l=0.05
R12 ui_in[5] a_24890_39160# sky130_fd_pr__res_generic_m2 w=0.45 l=0.05
X64 a_24200_41490# a_26090_39160# VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.35 pd=2.7 as=0.4 ps=2.8 w=1 l=0.15
X65 ua[0] a_23810_40680# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.189 pd=1.74 as=0.168 ps=1.64 w=0.42 l=0.15
X66 a_21880_39160# a_21880_39160# VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.35 pd=2.7 as=0.4 ps=2.8 w=1 l=0.15
X67 a_21880_39160# a_22770_39050# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.54 as=0.168 ps=1.64 w=0.42 l=0.15
X68 a_13100_38710# a_13070_38680# w_12870_38970# VGND sky130_fd_pr__nfet_01v8 ad=0.168 pd=1.64 as=0.189 ps=1.74 w=0.42 l=0.15
R13 uio_in[1] a_23250_39050# sky130_fd_pr__res_generic_m2 w=0.45 l=0.05
X69 a_21880_41750# a_21810_39050# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.54 as=0.168 ps=1.64 w=0.42 l=0.15
X70 a_24200_41490# a_24200_41490# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.54 as=0.168 ps=1.64 w=0.42 l=0.15
X71 ua[1] a_21880_39160# VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.55 pd=3.1 as=0.55 ps=3.1 w=1 l=0.15
X72 a_21880_41750# a_21880_41750# VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.35 pd=2.7 as=0.4 ps=2.8 w=1 l=0.15
X73 a_24200_41490# a_25610_39160# VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.35 pd=2.7 as=0.4 ps=2.8 w=1 l=0.15
X74 a_21880_39160# a_21880_39160# VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.35 pd=2.7 as=0.4 ps=2.8 w=1 l=0.15
X75 a_24200_38900# a_26090_39160# VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.35 pd=2.7 as=0.4 ps=2.8 w=1 l=0.15
X76 a_21880_39160# a_21810_39050# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.54 as=0.168 ps=1.64 w=0.42 l=0.15
X77 a_24200_38900# a_24200_38900# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.54 as=0.168 ps=1.64 w=0.42 l=0.15
R14 uio_in[7] a_21810_39050# sky130_fd_pr__res_generic_m2 w=0.45 l=0.05
R15 ui_in[1] a_25850_39160# sky130_fd_pr__res_generic_m2 w=0.45 l=0.05
C0 a_24890_39160# a_24200_41490# 0.220228f
C1 a_25130_39160# a_26090_39160# 1.13e-19
C2 a_25370_39160# a_25850_39160# 1.49e-19
C3 m2_22870_44110# uio_in[1] 0.021608f
C4 a_24650_39160# a_24200_41490# 0.219087f
C5 a_25130_39160# a_25850_39160# 1.34e-19
C6 a_25370_39160# a_25610_39160# 1.3709f
C7 a_24410_39160# a_24200_41490# 0.18266f
C8 a_24890_39160# a_25850_39160# 3.05e-19
C9 a_25130_39160# a_25610_39160# 1.56e-19
C10 m2_22130_44110# uio_in[2] 0.021608f
C11 a_24890_39160# a_25610_39160# 1.23e-19
C12 a_25130_39160# a_25370_39160# 1.31698f
C13 m2_28790_44110# m2_29530_44110# 0.007143f
C14 a_24890_39160# a_25370_39160# 1.78e-19
C15 m2_21390_44110# uio_in[3] 0.021608f
C16 a_24890_39160# a_25130_39160# 1.21119f
C17 m2_28050_44110# m2_28790_44110# 0.007143f
C18 a_24650_39160# a_25130_39160# 8.46e-19
C19 m2_20650_44110# uio_in[4] 0.021608f
C20 a_24650_39160# a_24890_39160# 1.10933f
C21 m2_27310_44110# m2_28050_44110# 0.007143f
C22 m2_19910_44110# uio_in[5] 0.021608f
C23 a_24410_39160# a_24650_39160# 1.01277f
C24 m2_26570_44110# m2_27310_44110# 0.007143f
C25 m2_19170_44110# uio_in[6] 0.021608f
C26 m2_25830_44110# m2_26570_44110# 0.007143f
C27 m2_18430_44110# uio_in[7] 0.021608f
C28 m2_25090_44110# m2_25830_44110# 0.007143f
C29 a_23490_39050# uio_in[0] 0.044617f
C30 a_26090_39160# ui_in[0] 0.049656f
C31 a_26090_39160# ui_in[1] 3.52e-19
C32 m2_24350_44110# m2_25090_44110# 0.007143f
C33 a_23250_39050# uio_in[1] 0.043751f
C34 a_25850_39160# ui_in[1] 0.049419f
C35 a_26090_39160# ui_in[2] 3.3e-19
C36 a_23010_39050# uio_in[1] 0.001582f
C37 a_25850_39160# ui_in[2] 5.76e-19
C38 a_26090_39160# ui_in[3] 3.3e-19
C39 a_23010_39050# uio_in[2] 0.046102f
C40 m2_23590_44110# m2_24350_44110# 0.006944f
C41 a_21880_41750# ua[1] 0.071522f
C42 a_24200_38900# ua[1] 0.023074f
C43 a_25850_39160# ui_in[3] 5.66e-19
C44 a_26090_39160# ui_in[4] 3.3e-19
C45 a_25610_39160# ui_in[2] 0.051252f
C46 a_22770_39050# uio_in[2] 0.001135f
C47 a_24200_38900# ua[0] 5.38e-20
C48 a_21880_39160# ua[1] 0.072223f
C49 a_25850_39160# ui_in[4] 5.53e-19
C50 a_25610_39160# ui_in[3] 6.72e-19
C51 a_22530_39050# uio_in[2] 8.23e-19
C52 a_22770_39050# uio_in[3] 0.047856f
C53 m2_22870_44110# m2_23590_44110# 0.007353f
C54 a_21880_41750# VPWR 1.67321f
C55 a_23810_40680# ua[1] 0.273365f
C56 a_25850_39160# ui_in[5] 0.001163f
C57 a_25370_39160# ui_in[3] 0.049254f
C58 a_25610_39160# ui_in[4] 6.57e-19
C59 a_24200_38900# VPWR 1.1585f
C60 a_22290_39050# uio_in[2] 6.38e-19
C61 a_22530_39050# uio_in[3] 8.23e-19
C62 a_23490_39050# ua[1] 0.092903f
C63 a_23810_40680# ua[0] 0.05951f
C64 a_25370_39160# ui_in[4] 8.82e-19
C65 a_25610_39160# ui_in[5] 6.45e-19
C66 a_21880_39160# VPWR 1.5973f
C67 a_22290_39050# uio_in[3] 6.38e-19
C68 a_22530_39050# uio_in[4] 0.049358f
C69 m2_22130_44110# m2_22870_44110# 0.007143f
C70 a_23250_39050# ua[1] 2.72e-19
C71 a_22050_39050# uio_in[3] 5.15e-19
C72 a_25130_39160# ui_in[4] 0.048012f
C73 a_25370_39160# ui_in[5] 8.67e-19
C74 a_23810_40680# VPWR 0.248173f
C75 a_22290_39050# uio_in[4] 6.38e-19
C76 a_23010_39050# ua[1] 1.47e-19
C77 a_21810_39050# uio_in[3] 2.96e-19
C78 a_22050_39050# uio_in[4] 5.15e-19
C79 a_25130_39160# ui_in[5] 0.001175f
C80 a_23490_39050# VPWR 0.534047f
C81 a_22290_39050# uio_in[5] 0.050403f
C82 m2_21390_44110# m2_22130_44110# 0.007143f
C83 a_22770_39050# ua[1] 9.1e-20
C84 a_21810_39050# uio_in[4] 2.96e-19
C85 a_22050_39050# uio_in[5] 5.15e-19
C86 a_24890_39160# ui_in[5] 0.046777f
C87 a_25130_39160# ui_in[6] 0.004014f
C88 a_23250_39050# VPWR 0.436562f
C89 m2_20650_44110# m2_21390_44110# 0.007143f
C90 a_22530_39050# ua[1] 6.16e-20
C91 a_21810_39050# uio_in[5] 2.96e-19
C92 a_22050_39050# uio_in[6] 0.051224f
C93 a_24890_39160# ui_in[6] 0.001608f
C94 a_23010_39050# VPWR 0.439864f
C95 a_22290_39050# ua[1] 4.44e-20
C96 a_21810_39050# uio_in[6] 2.96e-19
C97 a_24650_39160# ui_in[6] 0.044593f
C98 a_22770_39050# VPWR 0.445789f
C99 m2_19910_44110# m2_20650_44110# 0.007143f
C100 a_21810_39050# uio_in[7] 0.050442f
C101 a_22530_39050# VPWR 0.459327f
C102 clk ena 0.023797f
C103 a_24410_39160# ui_in[7] 0.044373f
C104 a_22290_39050# VPWR 0.478277f
C105 a_24200_41490# ua[1] 0.019982f
C106 m2_19170_44110# m2_19910_44110# 0.007143f
C107 a_22050_39050# VPWR 0.510229f
C108 rst_n clk 0.023797f
C109 a_26090_39160# ua[1] 1.8e-19
C110 a_24200_41490# ua[0] 0.001164f
C111 a_21810_39050# VPWR 0.87516f
C112 a_25850_39160# ua[1] 1.8e-19
C113 a_26090_39160# ua[0] 0.100513f
C114 m2_18430_44110# m2_19170_44110# 0.007143f
C115 a_24200_41490# VPWR 1.2358f
C116 ui_in[0] rst_n 0.023797f
C117 a_25850_39160# ua[0] 0.05653f
C118 a_25610_39160# ua[1] 1.8e-19
C119 a_26090_39160# VPWR 0.90977f
C120 a_25370_39160# ua[1] 1.8e-19
C121 a_25610_39160# ua[0] 0.055424f
C122 a_23490_39050# m2_23590_44110# 0.005112f
C123 a_25850_39160# VPWR 0.567946f
C124 ui_in[1] ui_in[0] 0.13387f
C125 a_26090_39160# m2_29530_44110# 0.005112f
C126 a_25130_39160# ua[1] 1.8e-19
C127 a_25370_39160# ua[0] 0.055026f
C128 a_25610_39160# VPWR 0.553411f
C129 li_14140_38880# m1_13270_38360# 0.057421f
C130 a_24890_39160# ua[1] 1.8e-19
C131 a_25130_39160# ua[0] 0.055076f
C132 a_23250_39050# m2_22870_44110# 0.005112f
C133 a_25370_39160# VPWR 0.537607f
C134 ui_in[2] ui_in[1] 0.133768f
C135 a_25130_39160# VPWR 0.527069f
C136 a_25850_39160# m2_28790_44110# 0.005112f
C137 a_13100_38710# m1_13270_38360# 0.0037f
C138 a_24650_39160# ua[1] 1.8e-19
C139 a_24890_39160# ua[0] 0.055733f
C140 a_24890_39160# VPWR 0.520247f
C141 a_13100_38710# li_14140_38880# 0.008859f
C142 a_24410_39160# ua[1] 0.093209f
C143 a_24650_39160# ua[0] 0.06855f
C144 a_23010_39050# m2_22130_44110# 0.005112f
C145 a_13070_38680# m1_13270_38360# 0.005568f
C146 ui_in[3] ui_in[2] 0.133458f
C147 a_24650_39160# VPWR 0.531904f
C148 a_25610_39160# m2_28050_44110# 0.005112f
C149 a_24410_39160# ua[0] 0.111655f
C150 a_13070_38680# li_14140_38880# 0.011142f
C151 w_12870_38970# m1_13270_38360# 0.00635f
C152 a_24410_39160# VPWR 0.663104f
C153 a_22770_39050# m2_21390_44110# 0.005112f
C154 a_13070_38680# a_13100_38710# 0.250071f
C155 w_12870_38970# li_14140_38880# 0.00761f
C156 ui_in[4] ui_in[3] 0.133435f
C157 a_25370_39160# m2_27310_44110# 0.005112f
C158 w_12870_38970# a_13100_38710# 0.411194f
C159 a_22530_39050# m2_20650_44110# 0.005112f
C160 w_12870_38970# a_13070_38680# 0.147772f
C161 ui_in[5] ui_in[4] 0.133252f
C162 a_25130_39160# m2_26570_44110# 0.005112f
C163 a_21880_39160# a_24200_38900# 0.001258f
C164 a_22290_39050# m2_19910_44110# 0.005112f
C165 a_21880_41750# a_23810_40680# 0.002387f
C166 ui_in[6] ui_in[5] 0.133228f
C167 a_23810_40680# a_24200_38900# 6.41e-21
C168 a_24890_39160# m2_25830_44110# 0.005112f
C169 a_21880_41750# a_23490_39050# 0.229552f
C170 a_23490_39050# a_24200_38900# 0.004679f
C171 a_23810_40680# a_21880_39160# 6.87e-19
C172 a_22050_39050# m2_19170_44110# 0.005112f
C173 a_21880_41750# a_23250_39050# 0.221622f
C174 ui_in[7] ui_in[6] 0.13321f
C175 a_23250_39050# a_24200_38900# 1.08e-20
C176 a_23490_39050# a_21880_39160# 0.21278f
C177 a_24650_39160# m2_25090_44110# 0.005112f
C178 a_21880_41750# a_23010_39050# 0.221772f
C179 VPWR ua[7] 0.010285f
C180 a_23010_39050# a_24200_38900# 6.92e-21
C181 a_23250_39050# a_21880_39160# 0.204846f
C182 a_23490_39050# a_23810_40680# 0.009378f
C183 a_21810_39050# m2_18430_44110# 0.005112f
C184 a_21880_41750# a_22770_39050# 0.222103f
C185 uio_in[0] ui_in[7] 0.132332f
C186 a_22770_39050# a_24200_38900# 4.79e-21
C187 a_23010_39050# a_21880_39160# 0.204812f
C188 a_23250_39050# a_23810_40680# 8.21e-19
C189 a_24410_39160# m2_24350_44110# 0.005112f
C190 a_21880_41750# a_22530_39050# 0.222316f
C191 a_22530_39050# a_24200_38900# 4.57e-22
C192 a_22770_39050# a_21880_39160# 0.204798f
C193 a_23010_39050# a_23810_40680# 4.18e-19
C194 a_23250_39050# a_23490_39050# 1.03051f
C195 a_21880_41750# a_22290_39050# 0.2225f
C196 uio_in[1] uio_in[0] 0.134137f
C197 a_22530_39050# a_21880_39160# 0.204791f
C198 a_22770_39050# a_23810_40680# 2.5e-19
C199 a_21880_41750# a_22050_39050# 0.222751f
C200 a_22290_39050# a_21880_39160# 0.204787f
C201 a_22530_39050# a_23810_40680# 1.65e-19
C202 a_23010_39050# a_23250_39050# 1.08328f
C203 a_21880_41750# a_21810_39050# 0.16944f
C204 uio_in[2] uio_in[1] 0.13321f
C205 a_22050_39050# a_21880_39160# 0.204778f
C206 a_22290_39050# a_23810_40680# 1.17e-19
C207 a_21880_41750# a_24200_41490# 0.001258f
C208 m2_29530_44110# ui_in[0] 0.020029f
C209 a_21810_39050# a_21880_39160# 0.159094f
C210 a_22770_39050# a_23010_39050# 1.19972f
C211 uio_in[3] uio_in[2] 0.13321f
C212 a_26090_39160# a_24200_38900# 0.143247f
C213 a_22530_39050# a_23010_39050# 1.6e-19
C214 m2_28790_44110# ui_in[1] 0.020255f
C215 VPWR ui_in[4] 0.004568f
C216 a_25850_39160# a_24200_38900# 0.143247f
C217 a_24200_41490# a_23810_40680# 0.001209f
C218 a_22290_39050# a_23010_39050# 1.13e-19
C219 a_22530_39050# a_22770_39050# 1.2778f
C220 uio_in[4] uio_in[3] 0.13321f
C221 VPWR ui_in[5] 0.004568f
C222 a_24200_41490# a_23490_39050# 0.004011f
C223 a_25610_39160# a_24200_38900# 0.143247f
C224 a_22290_39050# a_22770_39050# 1.23e-19
C225 a_21880_41750# a_25370_39160# 8.25e-21
C226 m2_28050_44110# ui_in[2] 0.02048f
C227 VPWR ui_in[6] 0.004568f
C228 a_24200_41490# a_23250_39050# 1.08e-20
C229 a_22050_39050# a_22770_39050# 9.52e-20
C230 a_25850_39160# a_23810_40680# 9.83e-20
C231 a_25370_39160# a_24200_38900# 0.143247f
C232 a_22290_39050# a_22530_39050# 1.45765f
C233 a_21880_41750# a_25130_39160# 1.16e-20
C234 uio_in[5] uio_in[4] 0.13321f
C235 VPWR ui_in[7] 0.004568f
C236 a_24200_41490# a_23010_39050# 6.92e-21
C237 a_22050_39050# a_22530_39050# 1.18e-19
C238 a_21810_39050# a_22770_39050# 7.47e-20
C239 a_25130_39160# a_24200_38900# 0.143247f
C240 a_25370_39160# a_21880_39160# 4.13e-21
C241 a_25610_39160# a_23810_40680# 1.39e-19
C242 a_21880_41750# a_24890_39160# 1.74e-20
C243 m2_27310_44110# ui_in[3] 0.020706f
C244 VPWR uio_in[0] 0.004568f
C245 a_24200_41490# a_22770_39050# 4.79e-21
C246 a_22050_39050# a_22290_39050# 1.64461f
C247 a_21810_39050# a_22530_39050# 9.71e-20
C248 a_24890_39160# a_24200_38900# 0.143247f
C249 a_25130_39160# a_21880_39160# 5.8e-21
C250 a_25370_39160# a_23810_40680# 2.12e-19
C251 a_21880_41750# a_24650_39160# 2.89e-20
C252 uio_in[6] uio_in[5] 0.13321f
C253 VPWR uio_in[1] 0.004568f
C254 a_24200_41490# a_22530_39050# 4.57e-22
C255 a_21810_39050# a_22290_39050# 1.06e-19
C256 a_24650_39160# a_24200_38900# 0.143247f
C257 a_24890_39160# a_21880_39160# 8.71e-21
C258 a_25130_39160# a_23810_40680# 3.6e-19
C259 a_21880_41750# a_24410_39160# 0.00727f
C260 VPWR uio_in[2] 0.004568f
C261 m2_26570_44110# ui_in[4] 0.020932f
C262 a_21810_39050# a_22050_39050# 1.66539f
C263 a_24410_39160# a_24200_38900# 0.111243f
C264 a_24650_39160# a_21880_39160# 1.44e-20
C265 a_24890_39160# a_23810_40680# 7.18e-19
C266 VPWR uio_in[3] 0.004568f
C267 uio_in[7] uio_in[6] 0.13321f
C268 a_24410_39160# a_21880_39160# 0.006714f
C269 a_24650_39160# a_23810_40680# 0.001837f
C270 VPWR uio_in[4] 0.004568f
C271 m2_25830_44110# ui_in[5] 0.021157f
C272 a_24410_39160# a_23810_40680# 0.049227f
C273 a_24410_39160# a_23490_39050# 0.222207f
C274 m2_25090_44110# ui_in[6] 0.021383f
C275 a_26090_39160# a_24200_41490# 0.215989f
C276 a_25850_39160# a_24200_41490# 0.221092f
C277 m2_24350_44110# ui_in[7] 0.021608f
C278 VPWR ua[1] 0.709125f
C279 a_25850_39160# a_26090_39160# 1.68469f
C280 a_25610_39160# a_24200_41490# 0.21981f
C281 VPWR ua[0] 0.765277f
C282 a_25370_39160# a_24200_41490# 0.220682f
C283 a_25610_39160# a_26090_39160# 1.54e-19
C284 m2_23590_44110# uio_in[0] 0.021608f
C285 a_25130_39160# a_24200_41490# 0.219289f
C286 a_25370_39160# a_26090_39160# 1.28e-19
C287 a_25610_39160# a_25850_39160# 1.89777f
C288 ua[2] VGND 0.122428f
C289 ua[3] VGND 0.122428f
C290 ua[4] VGND 0.122428f
C291 ua[5] VGND 0.122428f
C292 ua[6] VGND 0.122428f
C293 ua[7] VGND 0.111009f
C294 ena VGND 0.073297f
C295 clk VGND 0.0487f
C296 rst_n VGND 0.0487f
C297 ui_in[0] VGND 0.350951f
C298 ui_in[1] VGND 0.234234f
C299 ui_in[2] VGND 0.230502f
C300 ui_in[3] VGND 0.230704f
C301 ui_in[4] VGND 0.223397f
C302 ui_in[5] VGND 0.22191f
C303 ui_in[6] VGND 0.220814f
C304 ui_in[7] VGND 0.223871f
C305 uio_in[0] VGND 0.225466f
C306 uio_in[1] VGND 0.224179f
C307 uio_in[2] VGND 0.221286f
C308 uio_in[3] VGND 0.219592f
C309 uio_in[4] VGND 0.218871f
C310 uio_in[5] VGND 0.224716f
C311 uio_in[6] VGND 0.224366f
C312 uio_in[7] VGND 0.362103f
C313 ua[1] VGND 18.018312f
C314 ua[0] VGND 18.881802f
C315 VPWR VGND 64.375f
C316 m2_29530_44110# VGND 0.049454f $ **FLOATING
C317 m2_28790_44110# VGND 0.040694f $ **FLOATING
C318 m2_28050_44110# VGND 0.040694f $ **FLOATING
C319 m2_27310_44110# VGND 0.040694f $ **FLOATING
C320 m2_26570_44110# VGND 0.040694f $ **FLOATING
C321 m2_25830_44110# VGND 0.040694f $ **FLOATING
C322 m2_25090_44110# VGND 0.040694f $ **FLOATING
C323 m2_24350_44110# VGND 0.040877f $ **FLOATING
C324 m2_23590_44110# VGND 0.040687f $ **FLOATING
C325 m2_22870_44110# VGND 0.040504f $ **FLOATING
C326 m2_22130_44110# VGND 0.040694f $ **FLOATING
C327 m2_21390_44110# VGND 0.040694f $ **FLOATING
C328 m2_20650_44110# VGND 0.040694f $ **FLOATING
C329 m2_19910_44110# VGND 0.040694f $ **FLOATING
C330 m2_19170_44110# VGND 0.040694f $ **FLOATING
C331 m2_18430_44110# VGND 0.049454f $ **FLOATING
C332 m1_13270_38360# VGND 0.934988f $ **FLOATING
C333 li_14140_38880# VGND 0.665446f $ **FLOATING
C334 a_13100_38710# VGND 0.453185f
C335 a_13070_38680# VGND 0.542482f
C336 a_24200_38900# VGND 2.73692f
C337 a_21880_39160# VGND 1.994f
C338 a_23810_40680# VGND 0.712389f
C339 a_23490_39050# VGND 1.66046f
C340 a_23250_39050# VGND 1.41306f
C341 a_23010_39050# VGND 1.54891f
C342 a_22770_39050# VGND 1.64741f
C343 a_22530_39050# VGND 1.73515f
C344 a_22290_39050# VGND 1.80588f
C345 a_22050_39050# VGND 1.90533f
C346 a_21810_39050# VGND 3.17095f
C347 a_24200_41490# VGND 2.66092f
C348 a_26090_39160# VGND 2.90456f
C349 a_25850_39160# VGND 1.70481f
C350 a_25610_39160# VGND 1.62106f
C351 a_25370_39160# VGND 1.57552f
C352 a_25130_39160# VGND 1.47461f
C353 a_24890_39160# VGND 1.37037f
C354 a_24650_39160# VGND 1.22953f
C355 a_24410_39160# VGND 1.37675f
C356 a_21880_41750# VGND 1.92325f
C357 w_12870_38970# VGND 1.34935f


